VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO transmission_gate
  CLASS Core ;
  FOREIGN transmission_gate ;
  ORIGIN 0 0 ;
  SIZE 3.22 BY 2.72 ;
  SITE unithd ;
  PIN GN
    ANTENNAGATEAREA 0.082500 ;
    PORT
      LAYER li1 ;
        RECT 2.520 1.750 2.910 2.200 ;
    END
  END GN
  PIN G
    ANTENNAGATEAREA 0.082500 ;
    PORT
      LAYER li1 ;
        RECT 2.510 1.080 2.900 1.530 ;
    END
  END G
  PIN O
    ANTENNADIFFAREA 0.451000 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.600 2.220 2.100 ;
        RECT 1.980 0.940 2.190 1.600 ;
        RECT 1.870 0.640 2.220 0.940 ;
        RECT 2.410 0.640 2.800 0.910 ;
        RECT 1.870 0.440 2.800 0.640 ;
    END
  END O
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.530 0.290 2.380 1.100 ;
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.185 1.310 3.415 2.910 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.700 2.080 1.110 2.635 ;
        RECT 0.660 1.630 1.110 2.080 ;
        RECT 0.750 1.420 1.110 1.630 ;
        RECT 1.310 1.600 1.660 2.100 ;
        RECT 1.370 1.420 1.600 1.600 ;
        RECT 0.560 1.170 1.600 1.420 ;
        RECT 1.370 0.940 1.600 1.170 ;
        RECT 0.660 0.470 1.110 0.920 ;
        RECT 0.710 0.085 1.090 0.470 ;
        RECT 1.310 0.440 1.660 0.940 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
END transmission_gate
END LIBRARY

