.subckt CDC Reset Next_Edge_LowV Falling_Y Rising_Y Conversion_Finished V_LOW V_HIGH V_SENSE
X0 FALLING_COMP.INV_DM.O FALLING_COMP.SR_MEM.NANDQ.O V_GND V_GND V_LOW V_LOW FALLING_COMP.SR_MEM.NANDQb.O sky130_fd_sc_hd__nand2_1
X1 CLOCK_GEN.INV_R.O CLOCK_GEN.SR_Op.NANDQ.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.SR_Op.NANDQb.O sky130_fd_sc_hd__nand2_1
X2 FINISH_COMP.INV_DM.O FINISH_COMP.SR_MEM.NANDQ.O V_GND V_GND V_LOW V_LOW FINISH_COMP.SR_MEM.NANDQb.O sky130_fd_sc_hd__nand2_1
X3 CLOCK_GEN.NAND_DR.O CLOCK_GEN.SR_OE.NANDQ.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.SR_OE.NANDQb.O sky130_fd_sc_hd__nand2_1
X4 RISING_COMP.INV_DM.O RISING_COMP.SR_MEM.NANDQ.O V_GND V_GND V_LOW V_LOW RISING_COMP.SR_MEM.NANDQb.O sky130_fd_sc_hd__nand2_1
X5 FULL_COUNTER.COUNT_DFF.Q 1 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW CLOCK_GEN.NOT_CLK.O FULL_COUNTER.COUNT_DFF.Qb sky130_fd_sc_hd__dfbbn_1
X6 FULL_COUNTER.COUNT_DFF.Q V_GND V_GND V_LOW V_LOW 1 sky130_fd_sc_hd__inv_1
X7 2 V_GND V_GND V_LOW V_LOW 3 sky130_fd_sc_hd__inv_1
X8 4 V_GND V_GND V_LOW V_LOW 5 sky130_fd_sc_hd__inv_1
X9 6 V_GND V_GND V_LOW V_LOW 7 sky130_fd_sc_hd__inv_1
X10 8 V_GND V_GND V_LOW V_LOW 9 sky130_fd_sc_hd__inv_1
X11 10 V_GND V_GND V_LOW V_LOW 11 sky130_fd_sc_hd__inv_1
X12 12 V_GND V_GND V_LOW V_LOW 13 sky130_fd_sc_hd__inv_1
X13 14 V_GND V_GND V_LOW V_LOW 15 sky130_fd_sc_hd__inv_1
X14 16 V_GND V_GND V_LOW V_LOW 17 sky130_fd_sc_hd__inv_1
X15 18 V_GND V_GND V_LOW V_LOW 19 sky130_fd_sc_hd__inv_1
X16 20 V_GND V_GND V_LOW V_LOW 21 sky130_fd_sc_hd__inv_1
X17 22 V_GND V_GND V_LOW V_LOW 23 sky130_fd_sc_hd__inv_1
X18 24 V_GND V_GND V_LOW V_LOW 25 sky130_fd_sc_hd__inv_1
X19 26 V_GND V_GND V_LOW V_LOW 27 sky130_fd_sc_hd__inv_1
X20 28 V_GND V_GND V_LOW V_LOW 29 sky130_fd_sc_hd__inv_1
X21 30 V_GND V_GND V_LOW V_LOW 31 sky130_fd_sc_hd__inv_1
X22 32 V_GND V_GND V_LOW V_LOW 33 sky130_fd_sc_hd__inv_1
X23 34 V_GND V_GND V_LOW V_LOW 35 sky130_fd_sc_hd__inv_1
X24 36 V_GND V_GND V_LOW V_LOW 37 sky130_fd_sc_hd__inv_1
X25 38 V_GND V_GND V_LOW V_LOW 39 sky130_fd_sc_hd__inv_1
X26 2 3 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 1 40 sky130_fd_sc_hd__dfbbn_1
X27 4 5 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 3 41 sky130_fd_sc_hd__dfbbn_1
X28 6 7 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 5 42 sky130_fd_sc_hd__dfbbn_1
X29 8 9 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 7 43 sky130_fd_sc_hd__dfbbn_1
X30 10 11 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 9 44 sky130_fd_sc_hd__dfbbn_1
X31 12 13 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 11 45 sky130_fd_sc_hd__dfbbn_1
X32 14 15 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 13 46 sky130_fd_sc_hd__dfbbn_1
X33 16 17 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 15 47 sky130_fd_sc_hd__dfbbn_1
X34 18 19 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 17 48 sky130_fd_sc_hd__dfbbn_1
X35 20 21 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 19 49 sky130_fd_sc_hd__dfbbn_1
X36 22 23 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 21 50 sky130_fd_sc_hd__dfbbn_1
X37 24 25 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 23 51 sky130_fd_sc_hd__dfbbn_1
X38 26 27 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 25 52 sky130_fd_sc_hd__dfbbn_1
X39 28 29 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 27 53 sky130_fd_sc_hd__dfbbn_1
X40 30 31 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 29 54 sky130_fd_sc_hd__dfbbn_1
X41 32 33 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 31 55 sky130_fd_sc_hd__dfbbn_1
X42 34 35 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 33 56 sky130_fd_sc_hd__dfbbn_1
X43 36 37 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 35 57 sky130_fd_sc_hd__dfbbn_1
X44 38 39 FULL_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 37 58 sky130_fd_sc_hd__dfbbn_1
X45 RISING_COUNTER.COUNT_DFF.Q 59 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW RISING_COMP.NAND3_COMP.O RISING_COUNTER.COUNT_DFF.Qb sky130_fd_sc_hd__dfbbn_1
X46 RISING_COUNTER.COUNT_DFF.Q V_GND V_GND V_LOW V_LOW 59 sky130_fd_sc_hd__inv_1
X47 60 V_GND V_GND V_LOW V_LOW 61 sky130_fd_sc_hd__inv_1
X48 62 V_GND V_GND V_LOW V_LOW 63 sky130_fd_sc_hd__inv_1
X49 64 V_GND V_GND V_LOW V_LOW 65 sky130_fd_sc_hd__inv_1
X50 66 V_GND V_GND V_LOW V_LOW 67 sky130_fd_sc_hd__inv_1
X51 68 V_GND V_GND V_LOW V_LOW 69 sky130_fd_sc_hd__inv_1
X52 70 V_GND V_GND V_LOW V_LOW 71 sky130_fd_sc_hd__inv_1
X53 72 V_GND V_GND V_LOW V_LOW 73 sky130_fd_sc_hd__inv_1
X54 74 V_GND V_GND V_LOW V_LOW 75 sky130_fd_sc_hd__inv_1
X55 76 V_GND V_GND V_LOW V_LOW 77 sky130_fd_sc_hd__inv_1
X56 78 V_GND V_GND V_LOW V_LOW 79 sky130_fd_sc_hd__inv_1
X57 80 V_GND V_GND V_LOW V_LOW 81 sky130_fd_sc_hd__inv_1
X58 82 V_GND V_GND V_LOW V_LOW 83 sky130_fd_sc_hd__inv_1
X59 84 V_GND V_GND V_LOW V_LOW 85 sky130_fd_sc_hd__inv_1
X60 86 V_GND V_GND V_LOW V_LOW 87 sky130_fd_sc_hd__inv_1
X61 88 V_GND V_GND V_LOW V_LOW 89 sky130_fd_sc_hd__inv_1
X62 60 61 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 59 90 sky130_fd_sc_hd__dfbbn_1
X63 62 63 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 61 91 sky130_fd_sc_hd__dfbbn_1
X64 64 65 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 63 92 sky130_fd_sc_hd__dfbbn_1
X65 66 67 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 65 93 sky130_fd_sc_hd__dfbbn_1
X66 68 69 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 67 94 sky130_fd_sc_hd__dfbbn_1
X67 70 71 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 69 95 sky130_fd_sc_hd__dfbbn_1
X68 72 73 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 71 96 sky130_fd_sc_hd__dfbbn_1
X69 74 75 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 73 97 sky130_fd_sc_hd__dfbbn_1
X70 76 77 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 75 98 sky130_fd_sc_hd__dfbbn_1
X71 78 79 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 77 99 sky130_fd_sc_hd__dfbbn_1
X72 80 81 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 79 100 sky130_fd_sc_hd__dfbbn_1
X73 82 83 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 81 101 sky130_fd_sc_hd__dfbbn_1
X74 84 85 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 83 102 sky130_fd_sc_hd__dfbbn_1
X75 86 87 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 85 103 sky130_fd_sc_hd__dfbbn_1
X76 88 89 RISING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 87 104 sky130_fd_sc_hd__dfbbn_1
X77 FALLING_COUNTER.COUNT_DFF.Q 105 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW FALLING_COMP.NAND3_COMP.O FALLING_COUNTER.COUNT_DFF.Qb sky130_fd_sc_hd__dfbbn_1
X78 FALLING_COUNTER.COUNT_DFF.Q V_GND V_GND V_LOW V_LOW 105 sky130_fd_sc_hd__inv_1
X79 106 V_GND V_GND V_LOW V_LOW 107 sky130_fd_sc_hd__inv_1
X80 108 V_GND V_GND V_LOW V_LOW 109 sky130_fd_sc_hd__inv_1
X81 110 V_GND V_GND V_LOW V_LOW 111 sky130_fd_sc_hd__inv_1
X82 112 V_GND V_GND V_LOW V_LOW 113 sky130_fd_sc_hd__inv_1
X83 114 V_GND V_GND V_LOW V_LOW 115 sky130_fd_sc_hd__inv_1
X84 116 V_GND V_GND V_LOW V_LOW 117 sky130_fd_sc_hd__inv_1
X85 118 V_GND V_GND V_LOW V_LOW 119 sky130_fd_sc_hd__inv_1
X86 120 V_GND V_GND V_LOW V_LOW 121 sky130_fd_sc_hd__inv_1
X87 122 V_GND V_GND V_LOW V_LOW 123 sky130_fd_sc_hd__inv_1
X88 124 V_GND V_GND V_LOW V_LOW 125 sky130_fd_sc_hd__inv_1
X89 126 V_GND V_GND V_LOW V_LOW 127 sky130_fd_sc_hd__inv_1
X90 128 V_GND V_GND V_LOW V_LOW 129 sky130_fd_sc_hd__inv_1
X91 130 V_GND V_GND V_LOW V_LOW 131 sky130_fd_sc_hd__inv_1
X92 132 V_GND V_GND V_LOW V_LOW 133 sky130_fd_sc_hd__inv_1
X93 134 V_GND V_GND V_LOW V_LOW 135 sky130_fd_sc_hd__inv_1
X94 106 107 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 105 136 sky130_fd_sc_hd__dfbbn_1
X95 108 109 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 107 137 sky130_fd_sc_hd__dfbbn_1
X96 110 111 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 109 138 sky130_fd_sc_hd__dfbbn_1
X97 112 113 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 111 139 sky130_fd_sc_hd__dfbbn_1
X98 114 115 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 113 140 sky130_fd_sc_hd__dfbbn_1
X99 116 117 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 115 141 sky130_fd_sc_hd__dfbbn_1
X100 118 119 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 117 142 sky130_fd_sc_hd__dfbbn_1
X101 120 121 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 119 143 sky130_fd_sc_hd__dfbbn_1
X102 122 123 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 121 144 sky130_fd_sc_hd__dfbbn_1
X103 124 125 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 123 145 sky130_fd_sc_hd__dfbbn_1
X104 126 127 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 125 146 sky130_fd_sc_hd__dfbbn_1
X105 128 129 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 127 147 sky130_fd_sc_hd__dfbbn_1
X106 130 131 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 129 148 sky130_fd_sc_hd__dfbbn_1
X107 132 133 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 131 149 sky130_fd_sc_hd__dfbbn_1
X108 134 135 FALLING_COUNTER.RST_INV.O V_LOW V_GND V_GND V_LOW V_LOW 133 150 sky130_fd_sc_hd__dfbbn_1
X109 LOW_CHAIN.low_chain_inv16.O V_GND V_GND V_LOW V_LOW FALLING_COMP.INV_DM.O sky130_fd_sc_hd__inv_1
X110 FALLING_COMP.INV_DP.O FALLING_COMP.SR_MEM.NANDQb.O V_GND V_GND V_LOW V_LOW FALLING_COMP.SR_MEM.NANDQ.O sky130_fd_sc_hd__nand2_1
X111 FALLING_COMP.SR_MEM.NANDQ.O V_GND V_GND V_LOW V_LOW FALLING_COMP.INV_Q.O sky130_fd_sc_hd__inv_1
X112 FALLING_COMP.SR_MEM.NANDQb.O V_GND V_GND V_LOW V_LOW FALLING_COMP.INV_Qb.O sky130_fd_sc_hd__inv_1
X113 CAP_CHAIN.cap_chain_inv16.O LOW_CHAIN.low_chain_inv16.O V_GND V_GND V_LOW V_LOW FALLING_COMP.NAND2_COMP.O sky130_fd_sc_hd__nand2_1
X114 FALLING_COMP.INV_Qb.O FALLING_COMP.INV_DP.O FALLING_COMP.NAND3_COMP.O CLOCK_GEN.SR_OE.NANDQ.O sky130_fd_sc_hd__nand3_1
X115 FINISH_CHAIN.finish_chain_inv15.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.INV_F.O sky130_fd_sc_hd__inv_1
X116 FALLING_COMP.NAND2_COMP.O CLOCK_GEN.INV_F.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.NAND_DF.O sky130_fd_sc_hd__nand2_1
X117 CLOCK_GEN.NAND_DF.O CLOCK_GEN.SR_OE.NANDQb.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.SR_OE.NANDQ.O sky130_fd_sc_hd__nand2_1
X118 CLOCK_GEN.SR_OE.NANDQ.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.INV_OE.O sky130_fd_sc_hd__inv_1
X119 Reset V_GND V_GND V_LOW V_LOW CLOCK_GEN.INV_R.O sky130_fd_sc_hd__inv_1
X120 FINISH_COMP.NAND3_COMP.O CLOCK_GEN.SR_Op.NANDQb.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.SR_Op.NANDQ.O sky130_fd_sc_hd__nand2_1
X121 Reset CLOCK_GEN.SR_Op.NANDQ.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.NOR_CLK.O sky130_fd_sc_hd__nor2_1
X122 CLOCK_GEN.SR_OE.NANDQ.O CLOCK_GEN.NOR_CLK.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.NAND_CLK.O sky130_fd_sc_hd__nand2_1
X123 CLOCK_GEN.NAND_CLK.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.NOT_CLK.O sky130_fd_sc_hd__inv_1
X124 FINISH_CHAIN.finish_chain_inv16.O V_GND V_GND V_LOW V_LOW FINISH_COMP.INV_DM.O sky130_fd_sc_hd__inv_1
X125 FINISH_COMP.INV_DP.O FINISH_COMP.SR_MEM.NANDQb.O V_GND V_GND V_LOW V_LOW FINISH_COMP.SR_MEM.NANDQ.O sky130_fd_sc_hd__nand2_1
X126 FINISH_COMP.SR_MEM.NANDQ.O V_GND V_GND V_LOW V_LOW FINISH_COMP.INV_Q.O sky130_fd_sc_hd__inv_1
X127 FINISH_COMP.SR_MEM.NANDQb.O V_GND V_GND V_LOW V_LOW FINISH_COMP.INV_Qb.O sky130_fd_sc_hd__inv_1
X128 INV_RISING_CAP.O FINISH_CHAIN.finish_chain_inv16.O V_GND V_GND V_LOW V_LOW FINISH_COMP.NAND2_COMP.O sky130_fd_sc_hd__nand2_1
X129 FINISH_COMP.INV_Qb.O FINISH_COMP.INV_DP.O FINISH_COMP.NAND3_COMP.O CLOCK_GEN.INV_OE.O sky130_fd_sc_hd__nand3_1
X130 INV_RISING_LOW.O V_GND V_GND V_LOW V_LOW RISING_COMP.INV_DM.O sky130_fd_sc_hd__inv_1
X131 RISING_COMP.INV_DP.O RISING_COMP.SR_MEM.NANDQb.O V_GND V_GND V_LOW V_LOW RISING_COMP.SR_MEM.NANDQ.O sky130_fd_sc_hd__nand2_1
X132 RISING_COMP.SR_MEM.NANDQ.O V_GND V_GND V_LOW V_LOW RISING_COMP.INV_Q.O sky130_fd_sc_hd__inv_1
X133 RISING_COMP.SR_MEM.NANDQb.O V_GND V_GND V_LOW V_LOW RISING_COMP.INV_Qb.O sky130_fd_sc_hd__inv_1
X134 INV_RISING_CAP.O INV_RISING_LOW.O V_GND V_GND V_LOW V_LOW RISING_COMP.NAND2_COMP.O sky130_fd_sc_hd__nand2_1
X135 RISING_COMP.INV_Qb.O RISING_COMP.INV_DP.O RISING_COMP.NAND3_COMP.O CLOCK_GEN.INV_OE.O sky130_fd_sc_hd__nand3_1
X136 FINISH_CHAIN.finish_chain_inv1.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv2.O sky130_fd_sc_hd__inv_1
X137 FINISH_CHAIN.finish_chain_inv2.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv3.O sky130_fd_sc_hd__inv_1
X138 FINISH_CHAIN.finish_chain_inv3.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv4.O sky130_fd_sc_hd__inv_1
X139 FINISH_CHAIN.finish_chain_inv4.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv5.O sky130_fd_sc_hd__inv_1
X140 FINISH_CHAIN.finish_chain_inv5.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv6.O sky130_fd_sc_hd__inv_1
X141 FINISH_CHAIN.finish_chain_inv6.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv7.O sky130_fd_sc_hd__inv_1
X142 FINISH_CHAIN.finish_chain_inv7.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv8.O sky130_fd_sc_hd__inv_1
X143 FINISH_CHAIN.finish_chain_inv8.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv9.O sky130_fd_sc_hd__inv_1
X144 FINISH_CHAIN.finish_chain_inv9.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv10.O sky130_fd_sc_hd__inv_1
X145 FINISH_CHAIN.finish_chain_inv10.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv11.O sky130_fd_sc_hd__inv_1
X146 FINISH_CHAIN.finish_chain_inv11.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv12.O sky130_fd_sc_hd__inv_1
X147 FINISH_CHAIN.finish_chain_inv12.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv13.O sky130_fd_sc_hd__inv_1
X148 FINISH_CHAIN.finish_chain_inv13.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv14.O sky130_fd_sc_hd__inv_1
X149 FINISH_CHAIN.finish_chain_inv14.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv15.O sky130_fd_sc_hd__inv_1
X150 FINISH_CHAIN.finish_chain_inv15.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv16.O sky130_fd_sc_hd__inv_1
X151 CAP_CHAIN.cap_chain_inv1.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv2.O sky130_fd_sc_hd__inv_1
X152 CAP_CHAIN.cap_chain_inv2.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv3.O sky130_fd_sc_hd__inv_1
X153 CAP_CHAIN.cap_chain_inv3.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv4.O sky130_fd_sc_hd__inv_1
X154 CAP_CHAIN.cap_chain_inv4.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv5.O sky130_fd_sc_hd__inv_1
X155 CAP_CHAIN.cap_chain_inv5.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv6.O sky130_fd_sc_hd__inv_1
X156 CAP_CHAIN.cap_chain_inv6.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv7.O sky130_fd_sc_hd__inv_1
X157 CAP_CHAIN.cap_chain_inv7.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv8.O sky130_fd_sc_hd__inv_1
X158 CAP_CHAIN.cap_chain_inv8.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv9.O sky130_fd_sc_hd__inv_1
X159 CAP_CHAIN.cap_chain_inv9.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv10.O sky130_fd_sc_hd__inv_1
X160 CAP_CHAIN.cap_chain_inv10.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv11.O sky130_fd_sc_hd__inv_1
X161 CAP_CHAIN.cap_chain_inv11.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv12.O sky130_fd_sc_hd__inv_1
X162 CAP_CHAIN.cap_chain_inv12.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv13.O sky130_fd_sc_hd__inv_1
X163 CAP_CHAIN.cap_chain_inv13.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv14.O sky130_fd_sc_hd__inv_1
X164 CAP_CHAIN.cap_chain_inv14.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv15.O sky130_fd_sc_hd__inv_1
X165 CAP_CHAIN.cap_chain_inv15.O V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv16.O sky130_fd_sc_hd__inv_1
X166 LOW_CHAIN.low_chain_inv1.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv2.O sky130_fd_sc_hd__inv_1
X167 LOW_CHAIN.low_chain_inv2.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv3.O sky130_fd_sc_hd__inv_1
X168 LOW_CHAIN.low_chain_inv3.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv4.O sky130_fd_sc_hd__inv_1
X169 LOW_CHAIN.low_chain_inv4.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv5.O sky130_fd_sc_hd__inv_1
X170 LOW_CHAIN.low_chain_inv5.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv6.O sky130_fd_sc_hd__inv_1
X171 LOW_CHAIN.low_chain_inv6.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv7.O sky130_fd_sc_hd__inv_1
X172 LOW_CHAIN.low_chain_inv7.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv8.O sky130_fd_sc_hd__inv_1
X173 LOW_CHAIN.low_chain_inv8.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv9.O sky130_fd_sc_hd__inv_1
X174 LOW_CHAIN.low_chain_inv9.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv10.O sky130_fd_sc_hd__inv_1
X175 LOW_CHAIN.low_chain_inv10.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv11.O sky130_fd_sc_hd__inv_1
X176 LOW_CHAIN.low_chain_inv11.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv12.O sky130_fd_sc_hd__inv_1
X177 LOW_CHAIN.low_chain_inv12.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv13.O sky130_fd_sc_hd__inv_1
X178 LOW_CHAIN.low_chain_inv13.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv14.O sky130_fd_sc_hd__inv_1
X179 LOW_CHAIN.low_chain_inv14.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv15.O sky130_fd_sc_hd__inv_1
X180 LOW_CHAIN.low_chain_inv15.O V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv16.O sky130_fd_sc_hd__inv_1

X181 V_HIGH V_SENSE RESET V_HIGH V_GND transmission_gate

X182 V_GND V_HIGH V_GND INV_EDGE.O CLOCK_GEN.NOT_CLK.O V_HIGH Next_Edge_HighV SLC

X183 CLOCK_GEN.NOT_CLK.O V_GND V_GND V_LOW V_LOW INV_EDGE.O sky130_fd_sc_hd__inv_1
X184 Reset V_GND V_GND V_LOW V_LOW FULL_COUNTER.RST_INV.O sky130_fd_sc_hd__inv_1
X185 RISING_COMP.NAND2_COMP.O FINISH_CHAIN.finish_chain_inv15.O V_GND V_GND V_LOW V_LOW CLOCK_GEN.NAND_DR.O sky130_fd_sc_hd__nand2_1
X186 INV_RISING_CAP.O V_GND V_GND V_LOW V_LOW FINISH_COMP.INV_DP.O sky130_fd_sc_hd__inv_1
X187 Reset V_GND V_GND V_LOW V_LOW RISING_COUNTER.RST_INV.O sky130_fd_sc_hd__inv_1
X188 INV_RISING_CAP.O V_GND V_GND V_LOW V_LOW RISING_COMP.INV_DP.O sky130_fd_sc_hd__inv_1
X189 Reset V_GND V_GND V_LOW V_LOW FALLING_COUNTER.RST_INV.O sky130_fd_sc_hd__inv_1
X190 CAP_CHAIN.cap_chain_inv16.O V_GND V_GND V_LOW V_LOW FALLING_COMP.INV_DP.O sky130_fd_sc_hd__inv_1
X191 INV_RISING_LOW.O V_GND V_GND V_LOW V_LOW FINISH_CHAIN.finish_chain_inv1.O sky130_fd_sc_hd__inv_1
X192 CAP_CHAIN.cap_chain_inv16.O V_GND V_GND V_LOW V_LOW INV_RISING_CAP.O sky130_fd_sc_hd__inv_1
X193 LOW_CHAIN.low_chain_inv16.O V_GND V_GND V_LOW V_LOW INV_RISING_LOW.O sky130_fd_sc_hd__inv_1
X194 Next_Edge_HighV V_GND V_GND V_HIGH V_SENSE CAP_CHAIN.cap_chain_inv1.O sky130_fd_sc_hd__inv_1
X195 Next_Edge_HighV V_GND V_GND V_LOW V_LOW LOW_CHAIN.low_chain_inv1.O sky130_fd_sc_hd__inv_1
V0 Falling_Low LOW_CHAIN.O DC 0
V1 LOW_CHAIN.I Next_Edge_HighV DC 0
V2 Falling_Cap CAP_CHAIN.O DC 0
V3 CAP_CHAIN.I Next_Edge_HighV DC 0
V4 Rising_Low INV_RISING_LOW.O DC 0
V5 INV_RISING_LOW.I Falling_Low DC 0
V6 Rising_Cap INV_RISING_CAP.O DC 0
V7 INV_RISING_CAP.I Falling_Cap DC 0
V8 Finish_Low FINISH_CHAIN.O DC 0
V9 Finish_Delay FINISH_CHAIN.Ob DC 0
V10 FINISH_CHAIN.I Rising_Low DC 0
V11 Rising_Y RISING_COMP.Y DC 0
V12 Rising_Done RISING_COMP.Done DC 0
V13 RISING_COMP.Output_Enable Rising_Output_Enable DC 0
V14 RISING_COMP.D_Minus Rising_Low DC 0
V15 RISING_COMP.D_Plus Rising_Cap DC 0
V16 Finish FINISH_COMP.Y DC 0
V17 FINISH_COMP.Output_Enable Rising_Output_Enable DC 0
V18 FINISH_COMP.D_Minus Finish_Low DC 0
V19 FINISH_COMP.D_Plus Rising_Cap DC 0
V20 Conversion_Finished CLOCK_GEN.Conv_Finish DC 0
V21 Next_Edge_LowV CLOCK_GEN.Next_Edge DC 0
V22 Falling_Output_Enable CLOCK_GEN.OE_Falling DC 0
V23 Rising_Output_Enable CLOCK_GEN.OE_Rising DC 0
V24 CLOCK_GEN.Finish Finish DC 0
V25 CLOCK_GEN.Reset Reset DC 0
V26 CLOCK_GEN.Finish_Delay Finish_Delay DC 0
V27 CLOCK_GEN.Done_Falling Falling_Done DC 0
V28 CLOCK_GEN.Done_Rising Rising_Done DC 0
V29 Falling_Y FALLING_COMP.Y DC 0
V30 Falling_Done FALLING_COMP.Done DC 0
V31 FALLING_COMP.Output_Enable Falling_Output_Enable DC 0
V32 FALLING_COMP.D_Minus Falling_Low DC 0
V33 FALLING_COMP.D_Plus Falling_Cap DC 0
V34 D_SUB2.0 FALLING_COUNTER.O.0 DC 0
V35 D_SUB2.1 FALLING_COUNTER.O.1 DC 0
V36 D_SUB2.2 FALLING_COUNTER.O.2 DC 0
V37 D_SUB2.3 FALLING_COUNTER.O.3 DC 0
V38 D_SUB2.4 FALLING_COUNTER.O.4 DC 0
V39 D_SUB2.5 FALLING_COUNTER.O.5 DC 0
V40 D_SUB2.6 FALLING_COUNTER.O.6 DC 0
V41 D_SUB2.7 FALLING_COUNTER.O.7 DC 0
V42 D_SUB2.8 FALLING_COUNTER.O.8 DC 0
V43 D_SUB2.9 FALLING_COUNTER.O.9 DC 0
V44 D_SUB2.10 FALLING_COUNTER.O.10 DC 0
V45 D_SUB2.11 FALLING_COUNTER.O.11 DC 0
V46 D_SUB2.12 FALLING_COUNTER.O.12 DC 0
V47 D_SUB2.13 FALLING_COUNTER.O.13 DC 0
V48 D_SUB2.14 FALLING_COUNTER.O.14 DC 0
V49 D_SUB2.15 FALLING_COUNTER.O.15 DC 0
V50 FALLING_COUNTER.RST Reset DC 0
V51 FALLING_COUNTER.CLK Falling_Y DC 0
V52 D_SUB1.0 RISING_COUNTER.O.0 DC 0
V53 D_SUB1.1 RISING_COUNTER.O.1 DC 0
V54 D_SUB1.2 RISING_COUNTER.O.2 DC 0
V55 D_SUB1.3 RISING_COUNTER.O.3 DC 0
V56 D_SUB1.4 RISING_COUNTER.O.4 DC 0
V57 D_SUB1.5 RISING_COUNTER.O.5 DC 0
V58 D_SUB1.6 RISING_COUNTER.O.6 DC 0
V59 D_SUB1.7 RISING_COUNTER.O.7 DC 0
V60 D_SUB1.8 RISING_COUNTER.O.8 DC 0
V61 D_SUB1.9 RISING_COUNTER.O.9 DC 0
V62 D_SUB1.10 RISING_COUNTER.O.10 DC 0
V63 D_SUB1.11 RISING_COUNTER.O.11 DC 0
V64 D_SUB1.12 RISING_COUNTER.O.12 DC 0
V65 D_SUB1.13 RISING_COUNTER.O.13 DC 0
V66 D_SUB1.14 RISING_COUNTER.O.14 DC 0
V67 D_SUB1.15 RISING_COUNTER.O.15 DC 0
V68 RISING_COUNTER.RST Reset DC 0
V69 RISING_COUNTER.CLK Rising_Y DC 0
V70 D_MAIN.0 FULL_COUNTER.O.0 DC 0
V71 D_MAIN.1 FULL_COUNTER.O.1 DC 0
V72 D_MAIN.2 FULL_COUNTER.O.2 DC 0
V73 D_MAIN.3 FULL_COUNTER.O.3 DC 0
V74 D_MAIN.4 FULL_COUNTER.O.4 DC 0
V75 D_MAIN.5 FULL_COUNTER.O.5 DC 0
V76 D_MAIN.6 FULL_COUNTER.O.6 DC 0
V77 D_MAIN.7 FULL_COUNTER.O.7 DC 0
V78 D_MAIN.8 FULL_COUNTER.O.8 DC 0
V79 D_MAIN.9 FULL_COUNTER.O.9 DC 0
V80 D_MAIN.10 FULL_COUNTER.O.10 DC 0
V81 D_MAIN.11 FULL_COUNTER.O.11 DC 0
V82 D_MAIN.12 FULL_COUNTER.O.12 DC 0
V83 D_MAIN.13 FULL_COUNTER.O.13 DC 0
V84 D_MAIN.14 FULL_COUNTER.O.14 DC 0
V85 D_MAIN.15 FULL_COUNTER.O.15 DC 0
V86 D_MAIN.16 FULL_COUNTER.O.16 DC 0
V87 D_MAIN.17 FULL_COUNTER.O.17 DC 0
V88 D_MAIN.18 FULL_COUNTER.O.18 DC 0
V89 D_MAIN.19 FULL_COUNTER.O.19 DC 0
V90 FULL_COUNTER.RST Reset DC 0
V91 FULL_COUNTER.CLK Next_Edge_LowV DC 0
V92 Next_Edge_LowV_b INV_EDGE.O DC 0
V93 INV_EDGE.I Next_Edge_LowV DC 0
V94 LOW_CHAIN.low_chain1 LOW_CHAIN.low_chain_inv1.O DC 0
V95 LOW_CHAIN.low_chain_inv1.I LOW_CHAIN.I DC 0
V96 LOW_CHAIN.low_chain2 LOW_CHAIN.low_chain_inv2.O DC 0
V97 LOW_CHAIN.low_chain_inv2.I LOW_CHAIN.low_chain1 DC 0
V98 LOW_CHAIN.low_chain3 LOW_CHAIN.low_chain_inv3.O DC 0
V99 LOW_CHAIN.low_chain_inv3.I LOW_CHAIN.low_chain2 DC 0
V100 LOW_CHAIN.low_chain4 LOW_CHAIN.low_chain_inv4.O DC 0
V101 LOW_CHAIN.low_chain_inv4.I LOW_CHAIN.low_chain3 DC 0
V102 LOW_CHAIN.low_chain5 LOW_CHAIN.low_chain_inv5.O DC 0
V103 LOW_CHAIN.low_chain_inv5.I LOW_CHAIN.low_chain4 DC 0
V104 LOW_CHAIN.low_chain6 LOW_CHAIN.low_chain_inv6.O DC 0
V105 LOW_CHAIN.low_chain_inv6.I LOW_CHAIN.low_chain5 DC 0
V106 LOW_CHAIN.low_chain7 LOW_CHAIN.low_chain_inv7.O DC 0
V107 LOW_CHAIN.low_chain_inv7.I LOW_CHAIN.low_chain6 DC 0
V108 LOW_CHAIN.low_chain8 LOW_CHAIN.low_chain_inv8.O DC 0
V109 LOW_CHAIN.low_chain_inv8.I LOW_CHAIN.low_chain7 DC 0
V110 LOW_CHAIN.low_chain9 LOW_CHAIN.low_chain_inv9.O DC 0
V111 LOW_CHAIN.low_chain_inv9.I LOW_CHAIN.low_chain8 DC 0
V112 LOW_CHAIN.low_chain10 LOW_CHAIN.low_chain_inv10.O DC 0
V113 LOW_CHAIN.low_chain_inv10.I LOW_CHAIN.low_chain9 DC 0
V114 LOW_CHAIN.low_chain11 LOW_CHAIN.low_chain_inv11.O DC 0
V115 LOW_CHAIN.low_chain_inv11.I LOW_CHAIN.low_chain10 DC 0
V116 LOW_CHAIN.low_chain12 LOW_CHAIN.low_chain_inv12.O DC 0
V117 LOW_CHAIN.low_chain_inv12.I LOW_CHAIN.low_chain11 DC 0
V118 LOW_CHAIN.low_chain13 LOW_CHAIN.low_chain_inv13.O DC 0
V119 LOW_CHAIN.low_chain_inv13.I LOW_CHAIN.low_chain12 DC 0
V120 LOW_CHAIN.low_chain14 LOW_CHAIN.low_chain_inv14.O DC 0
V121 LOW_CHAIN.low_chain_inv14.I LOW_CHAIN.low_chain13 DC 0
V122 LOW_CHAIN.low_chain15 LOW_CHAIN.low_chain_inv15.O DC 0
V123 LOW_CHAIN.low_chain_inv15.I LOW_CHAIN.low_chain14 DC 0
V124 LOW_CHAIN.O LOW_CHAIN.low_chain_inv16.O DC 0
V125 LOW_CHAIN.low_chain_inv16.I LOW_CHAIN.low_chain15 DC 0
V126 CAP_CHAIN.cap_chain1 CAP_CHAIN.cap_chain_inv1.O DC 0
V127 CAP_CHAIN.cap_chain_inv1.I CAP_CHAIN.I DC 0
V128 CAP_CHAIN.cap_chain2 CAP_CHAIN.cap_chain_inv2.O DC 0
V129 CAP_CHAIN.cap_chain_inv2.I CAP_CHAIN.cap_chain1 DC 0
V130 CAP_CHAIN.cap_chain3 CAP_CHAIN.cap_chain_inv3.O DC 0
V131 CAP_CHAIN.cap_chain_inv3.I CAP_CHAIN.cap_chain2 DC 0
V132 CAP_CHAIN.cap_chain4 CAP_CHAIN.cap_chain_inv4.O DC 0
V133 CAP_CHAIN.cap_chain_inv4.I CAP_CHAIN.cap_chain3 DC 0
V134 CAP_CHAIN.cap_chain5 CAP_CHAIN.cap_chain_inv5.O DC 0
V135 CAP_CHAIN.cap_chain_inv5.I CAP_CHAIN.cap_chain4 DC 0
V136 CAP_CHAIN.cap_chain6 CAP_CHAIN.cap_chain_inv6.O DC 0
V137 CAP_CHAIN.cap_chain_inv6.I CAP_CHAIN.cap_chain5 DC 0
V138 CAP_CHAIN.cap_chain7 CAP_CHAIN.cap_chain_inv7.O DC 0
V139 CAP_CHAIN.cap_chain_inv7.I CAP_CHAIN.cap_chain6 DC 0
V140 CAP_CHAIN.cap_chain8 CAP_CHAIN.cap_chain_inv8.O DC 0
V141 CAP_CHAIN.cap_chain_inv8.I CAP_CHAIN.cap_chain7 DC 0
V142 CAP_CHAIN.cap_chain9 CAP_CHAIN.cap_chain_inv9.O DC 0
V143 CAP_CHAIN.cap_chain_inv9.I CAP_CHAIN.cap_chain8 DC 0
V144 CAP_CHAIN.cap_chain10 CAP_CHAIN.cap_chain_inv10.O DC 0
V145 CAP_CHAIN.cap_chain_inv10.I CAP_CHAIN.cap_chain9 DC 0
V146 CAP_CHAIN.cap_chain11 CAP_CHAIN.cap_chain_inv11.O DC 0
V147 CAP_CHAIN.cap_chain_inv11.I CAP_CHAIN.cap_chain10 DC 0
V148 CAP_CHAIN.cap_chain12 CAP_CHAIN.cap_chain_inv12.O DC 0
V149 CAP_CHAIN.cap_chain_inv12.I CAP_CHAIN.cap_chain11 DC 0
V150 CAP_CHAIN.cap_chain13 CAP_CHAIN.cap_chain_inv13.O DC 0
V151 CAP_CHAIN.cap_chain_inv13.I CAP_CHAIN.cap_chain12 DC 0
V152 CAP_CHAIN.cap_chain14 CAP_CHAIN.cap_chain_inv14.O DC 0
V153 CAP_CHAIN.cap_chain_inv14.I CAP_CHAIN.cap_chain13 DC 0
V154 CAP_CHAIN.cap_chain15 CAP_CHAIN.cap_chain_inv15.O DC 0
V155 CAP_CHAIN.cap_chain_inv15.I CAP_CHAIN.cap_chain14 DC 0
V156 CAP_CHAIN.O CAP_CHAIN.cap_chain_inv16.O DC 0
V157 CAP_CHAIN.cap_chain_inv16.I CAP_CHAIN.cap_chain15 DC 0
V158 FINISH_CHAIN.finish_chain1 FINISH_CHAIN.finish_chain_inv1.O DC 0
V159 FINISH_CHAIN.finish_chain_inv1.I FINISH_CHAIN.I DC 0
V160 FINISH_CHAIN.finish_chain2 FINISH_CHAIN.finish_chain_inv2.O DC 0
V161 FINISH_CHAIN.finish_chain_inv2.I FINISH_CHAIN.finish_chain1 DC 0
V162 FINISH_CHAIN.finish_chain3 FINISH_CHAIN.finish_chain_inv3.O DC 0
V163 FINISH_CHAIN.finish_chain_inv3.I FINISH_CHAIN.finish_chain2 DC 0
V164 FINISH_CHAIN.finish_chain4 FINISH_CHAIN.finish_chain_inv4.O DC 0
V165 FINISH_CHAIN.finish_chain_inv4.I FINISH_CHAIN.finish_chain3 DC 0
V166 FINISH_CHAIN.finish_chain5 FINISH_CHAIN.finish_chain_inv5.O DC 0
V167 FINISH_CHAIN.finish_chain_inv5.I FINISH_CHAIN.finish_chain4 DC 0
V168 FINISH_CHAIN.finish_chain6 FINISH_CHAIN.finish_chain_inv6.O DC 0
V169 FINISH_CHAIN.finish_chain_inv6.I FINISH_CHAIN.finish_chain5 DC 0
V170 FINISH_CHAIN.finish_chain7 FINISH_CHAIN.finish_chain_inv7.O DC 0
V171 FINISH_CHAIN.finish_chain_inv7.I FINISH_CHAIN.finish_chain6 DC 0
V172 FINISH_CHAIN.finish_chain8 FINISH_CHAIN.finish_chain_inv8.O DC 0
V173 FINISH_CHAIN.finish_chain_inv8.I FINISH_CHAIN.finish_chain7 DC 0
V174 FINISH_CHAIN.finish_chain9 FINISH_CHAIN.finish_chain_inv9.O DC 0
V175 FINISH_CHAIN.finish_chain_inv9.I FINISH_CHAIN.finish_chain8 DC 0
V176 FINISH_CHAIN.finish_chain10 FINISH_CHAIN.finish_chain_inv10.O DC 0
V177 FINISH_CHAIN.finish_chain_inv10.I FINISH_CHAIN.finish_chain9 DC 0
V178 FINISH_CHAIN.finish_chain11 FINISH_CHAIN.finish_chain_inv11.O DC 0
V179 FINISH_CHAIN.finish_chain_inv11.I FINISH_CHAIN.finish_chain10 DC 0
V180 FINISH_CHAIN.finish_chain12 FINISH_CHAIN.finish_chain_inv12.O DC 0
V181 FINISH_CHAIN.finish_chain_inv12.I FINISH_CHAIN.finish_chain11 DC 0
V182 FINISH_CHAIN.finish_chain13 FINISH_CHAIN.finish_chain_inv13.O DC 0
V183 FINISH_CHAIN.finish_chain_inv13.I FINISH_CHAIN.finish_chain12 DC 0
V184 FINISH_CHAIN.finish_chain14 FINISH_CHAIN.finish_chain_inv14.O DC 0
V185 FINISH_CHAIN.finish_chain_inv14.I FINISH_CHAIN.finish_chain13 DC 0
V186 FINISH_CHAIN.Ob FINISH_CHAIN.finish_chain_inv15.O DC 0
V187 FINISH_CHAIN.finish_chain_inv15.I FINISH_CHAIN.finish_chain14 DC 0
V188 FINISH_CHAIN.O FINISH_CHAIN.finish_chain_inv16.O DC 0
V189 FINISH_CHAIN.finish_chain_inv16.I FINISH_CHAIN.Ob DC 0
V190 RISING_COMP.Db_Minus RISING_COMP.INV_DM.O DC 0
V191 RISING_COMP.INV_DM.I RISING_COMP.D_Minus DC 0
V192 RISING_COMP.Db_Plus RISING_COMP.INV_DP.O DC 0
V193 RISING_COMP.INV_DP.I RISING_COMP.D_Plus DC 0
V194 RISING_COMP.Qb RISING_COMP.SR_MEM.Qb DC 0
V195 RISING_COMP.Q RISING_COMP.SR_MEM.Q DC 0
V196 RISING_COMP.SR_MEM.Rb RISING_COMP.Db_Minus DC 0
V197 RISING_COMP.SR_MEM.Sb RISING_COMP.Db_Plus DC 0
V198 RISING_COMP.Qb_b RISING_COMP.INV_Qb.O DC 0
V199 RISING_COMP.INV_Qb.I RISING_COMP.Qb DC 0
V200 CLOCK_GEN.FinishB_Delay CLOCK_GEN.INV_F.O DC 0
V201 CLOCK_GEN.INV_F.I CLOCK_GEN.Finish_Delay DC 0
V202 FALLING_COMP.Done FALLING_COMP.NAND2_COMP.O DC 0
V203 FALLING_COMP.NAND2_COMP.B FALLING_COMP.D_Minus DC 0
V204 FALLING_COMP.NAND2_COMP.A FALLING_COMP.D_Plus DC 0
V205 CLOCK_GEN.Set_OE CLOCK_GEN.NAND_DF.O DC 0
V206 CLOCK_GEN.NAND_DF.B CLOCK_GEN.FinishB_Delay DC 0
V207 CLOCK_GEN.NAND_DF.A CLOCK_GEN.Done_Falling DC 0
V208 RISING_COMP.Done RISING_COMP.NAND2_COMP.O DC 0
V209 RISING_COMP.NAND2_COMP.B RISING_COMP.D_Minus DC 0
V210 RISING_COMP.NAND2_COMP.A RISING_COMP.D_Plus DC 0
V211 CLOCK_GEN.Reset_OE CLOCK_GEN.NAND_DR.O DC 0
V212 CLOCK_GEN.NAND_DR.B CLOCK_GEN.Finish_Delay DC 0
V213 CLOCK_GEN.NAND_DR.A CLOCK_GEN.Done_Rising DC 0
V214 CLOCK_GEN.OE_Falling CLOCK_GEN.SR_OE.Q DC 0
V215 CLOCK_GEN.SR_OE.Rb CLOCK_GEN.Reset_OE DC 0
V216 CLOCK_GEN.SR_OE.Sb CLOCK_GEN.Set_OE DC 0
V217 CLOCK_GEN.OE_Rising CLOCK_GEN.INV_OE.O DC 0
V218 CLOCK_GEN.INV_OE.I CLOCK_GEN.OE_Falling DC 0
V219 RISING_COMP.Y RISING_COMP.NAND3_COMP.O DC 0
V220 RISING_COMP.NAND3_COMP.C RISING_COMP.Output_Enable DC 0
V221 RISING_COMP.NAND3_COMP.B RISING_COMP.Db_Plus DC 0
V222 RISING_COMP.NAND3_COMP.A RISING_COMP.Qb_b DC 0
V223 RISING_COMP.Q_b RISING_COMP.INV_Q.O DC 0
V224 RISING_COMP.INV_Q.I RISING_COMP.Q DC 0
V225 FINISH_COMP.Db_Minus FINISH_COMP.INV_DM.O DC 0
V226 FINISH_COMP.INV_DM.I FINISH_COMP.D_Minus DC 0
V227 FINISH_COMP.Db_Plus FINISH_COMP.INV_DP.O DC 0
V228 FINISH_COMP.INV_DP.I FINISH_COMP.D_Plus DC 0
V229 FINISH_COMP.Qb FINISH_COMP.SR_MEM.Qb DC 0
V230 FINISH_COMP.Q FINISH_COMP.SR_MEM.Q DC 0
V231 FINISH_COMP.SR_MEM.Rb FINISH_COMP.Db_Minus DC 0
V232 FINISH_COMP.SR_MEM.Sb FINISH_COMP.Db_Plus DC 0
V233 FINISH_COMP.Qb_b FINISH_COMP.INV_Qb.O DC 0
V234 FINISH_COMP.INV_Qb.I FINISH_COMP.Qb DC 0
V235 FINISH_COMP.Y FINISH_COMP.NAND3_COMP.O DC 0
V236 FINISH_COMP.NAND3_COMP.C FINISH_COMP.Output_Enable DC 0
V237 FINISH_COMP.NAND3_COMP.B FINISH_COMP.Db_Plus DC 0
V238 FINISH_COMP.NAND3_COMP.A FINISH_COMP.Qb_b DC 0
V239 FINISH_COMP.Done FINISH_COMP.NAND2_COMP.O DC 0
V240 FINISH_COMP.NAND2_COMP.B FINISH_COMP.D_Minus DC 0
V241 FINISH_COMP.NAND2_COMP.A FINISH_COMP.D_Plus DC 0
V242 FINISH_COMP.Q_b FINISH_COMP.INV_Q.O DC 0
V243 FINISH_COMP.INV_Q.I FINISH_COMP.Q DC 0
V244 CLOCK_GEN.ResetB CLOCK_GEN.INV_R.O DC 0
V245 CLOCK_GEN.INV_R.I CLOCK_GEN.Reset DC 0
V246 CLOCK_GEN.Conv_Finish CLOCK_GEN.SR_Op.Q DC 0
V247 CLOCK_GEN.SR_Op.Rb CLOCK_GEN.ResetB DC 0
V248 CLOCK_GEN.SR_Op.Sb CLOCK_GEN.Finish DC 0
V249 CLOCK_GEN.Sense CLOCK_GEN.NOR_CLK.O DC 0
V250 CLOCK_GEN.NOR_CLK.B CLOCK_GEN.Conv_Finish DC 0
V251 CLOCK_GEN.NOR_CLK.A CLOCK_GEN.Reset DC 0
V252 CLOCK_GEN.CLKb CLOCK_GEN.NAND_CLK.O DC 0
V253 CLOCK_GEN.NAND_CLK.B CLOCK_GEN.Sense DC 0
V254 CLOCK_GEN.NAND_CLK.A CLOCK_GEN.OE_Falling DC 0
V255 CLOCK_GEN.Next_Edge CLOCK_GEN.NOT_CLK.O DC 0
V256 CLOCK_GEN.NOT_CLK.I CLOCK_GEN.CLKb DC 0
V257 FALLING_COMP.Db_Minus FALLING_COMP.INV_DM.O DC 0
V258 FALLING_COMP.INV_DM.I FALLING_COMP.D_Minus DC 0
V259 FALLING_COMP.Db_Plus FALLING_COMP.INV_DP.O DC 0
V260 FALLING_COMP.INV_DP.I FALLING_COMP.D_Plus DC 0
V261 FALLING_COMP.Qb FALLING_COMP.SR_MEM.Qb DC 0
V262 FALLING_COMP.Q FALLING_COMP.SR_MEM.Q DC 0
V263 FALLING_COMP.SR_MEM.Rb FALLING_COMP.Db_Minus DC 0
V264 FALLING_COMP.SR_MEM.Sb FALLING_COMP.Db_Plus DC 0
V265 FALLING_COMP.Qb_b FALLING_COMP.INV_Qb.O DC 0
V266 FALLING_COMP.INV_Qb.I FALLING_COMP.Qb DC 0
V267 FALLING_COUNTER.D.14 133 DC 0
V268 151 FALLING_COUNTER.O.14 DC 0
V269 FALLING_COMP.Y FALLING_COMP.NAND3_COMP.O DC 0
V270 FALLING_COMP.NAND3_COMP.C FALLING_COMP.Output_Enable DC 0
V271 FALLING_COMP.NAND3_COMP.B FALLING_COMP.Db_Plus DC 0
V272 FALLING_COMP.NAND3_COMP.A FALLING_COMP.Qb_b DC 0
V273 FALLING_COUNTER.RSTb FALLING_COUNTER.RST_INV.O DC 0
V274 FALLING_COUNTER.RST_INV.I FALLING_COUNTER.RST DC 0
V275 FALLING_COUNTER.O.0 FALLING_COUNTER.COUNT_DFF.Q DC 0
V276 FALLING_COUNTER.COUNT_DFF.RSTb FALLING_COUNTER.RSTb DC 0
V277 FALLING_COUNTER.COUNT_DFF.D FALLING_COUNTER.D.0 DC 0
V278 FALLING_COUNTER.COUNT_DFF.CLK FALLING_COUNTER.CLK DC 0
V279 FALLING_COUNTER.D.0 105 DC 0
V280 152 FALLING_COUNTER.O.0 DC 0
V281 FALLING_COUNTER.O.1 106 DC 0
V282 153 FALLING_COUNTER.RSTb DC 0
V283 154 FALLING_COUNTER.D.1 DC 0
V284 155 FALLING_COUNTER.D.0 DC 0
V285 FALLING_COUNTER.D.1 107 DC 0
V286 156 FALLING_COUNTER.O.1 DC 0
V287 FALLING_COUNTER.O.2 108 DC 0
V288 157 FALLING_COUNTER.RSTb DC 0
V289 158 FALLING_COUNTER.D.2 DC 0
V290 159 FALLING_COUNTER.D.1 DC 0
V291 FALLING_COUNTER.D.2 109 DC 0
V292 160 FALLING_COUNTER.O.2 DC 0
V293 FALLING_COUNTER.O.3 110 DC 0
V294 161 FALLING_COUNTER.RSTb DC 0
V295 162 FALLING_COUNTER.D.3 DC 0
V296 163 FALLING_COUNTER.D.2 DC 0
V297 FALLING_COUNTER.D.3 111 DC 0
V298 164 FALLING_COUNTER.O.3 DC 0
V299 FALLING_COUNTER.O.4 112 DC 0
V300 165 FALLING_COUNTER.RSTb DC 0
V301 166 FALLING_COUNTER.D.4 DC 0
V302 167 FALLING_COUNTER.D.3 DC 0
V303 FALLING_COUNTER.D.4 113 DC 0
V304 168 FALLING_COUNTER.O.4 DC 0
V305 FALLING_COUNTER.O.5 114 DC 0
V306 169 FALLING_COUNTER.RSTb DC 0
V307 170 FALLING_COUNTER.D.5 DC 0
V308 171 FALLING_COUNTER.D.4 DC 0
V309 FALLING_COUNTER.D.5 115 DC 0
V310 172 FALLING_COUNTER.O.5 DC 0
V311 FALLING_COUNTER.O.6 116 DC 0
V312 173 FALLING_COUNTER.RSTb DC 0
V313 174 FALLING_COUNTER.D.6 DC 0
V314 175 FALLING_COUNTER.D.5 DC 0
V315 FALLING_COUNTER.D.6 117 DC 0
V316 176 FALLING_COUNTER.O.6 DC 0
V317 FALLING_COUNTER.O.7 118 DC 0
V318 177 FALLING_COUNTER.RSTb DC 0
V319 178 FALLING_COUNTER.D.7 DC 0
V320 179 FALLING_COUNTER.D.6 DC 0
V321 FALLING_COUNTER.D.7 119 DC 0
V322 180 FALLING_COUNTER.O.7 DC 0
V323 FALLING_COUNTER.O.8 120 DC 0
V324 181 FALLING_COUNTER.RSTb DC 0
V325 182 FALLING_COUNTER.D.8 DC 0
V326 183 FALLING_COUNTER.D.7 DC 0
V327 FALLING_COUNTER.D.8 121 DC 0
V328 184 FALLING_COUNTER.O.8 DC 0
V329 FALLING_COUNTER.O.9 122 DC 0
V330 185 FALLING_COUNTER.RSTb DC 0
V331 186 FALLING_COUNTER.D.9 DC 0
V332 187 FALLING_COUNTER.D.8 DC 0
V333 FALLING_COUNTER.D.9 123 DC 0
V334 188 FALLING_COUNTER.O.9 DC 0
V335 FALLING_COUNTER.O.10 124 DC 0
V336 189 FALLING_COUNTER.RSTb DC 0
V337 190 FALLING_COUNTER.D.10 DC 0
V338 191 FALLING_COUNTER.D.9 DC 0
V339 FALLING_COUNTER.D.10 125 DC 0
V340 192 FALLING_COUNTER.O.10 DC 0
V341 FALLING_COUNTER.O.11 126 DC 0
V342 193 FALLING_COUNTER.RSTb DC 0
V343 194 FALLING_COUNTER.D.11 DC 0
V344 195 FALLING_COUNTER.D.10 DC 0
V345 FALLING_COUNTER.D.11 127 DC 0
V346 196 FALLING_COUNTER.O.11 DC 0
V347 FALLING_COUNTER.O.12 128 DC 0
V348 197 FALLING_COUNTER.RSTb DC 0
V349 198 FALLING_COUNTER.D.12 DC 0
V350 199 FALLING_COUNTER.D.11 DC 0
V351 FALLING_COUNTER.D.12 129 DC 0
V352 200 FALLING_COUNTER.O.12 DC 0
V353 FALLING_COUNTER.O.13 130 DC 0
V354 201 FALLING_COUNTER.RSTb DC 0
V355 202 FALLING_COUNTER.D.13 DC 0
V356 203 FALLING_COUNTER.D.12 DC 0
V357 FALLING_COUNTER.D.13 131 DC 0
V358 204 FALLING_COUNTER.O.13 DC 0
V359 FALLING_COUNTER.O.14 132 DC 0
V360 205 FALLING_COUNTER.RSTb DC 0
V361 206 FALLING_COUNTER.D.14 DC 0
V362 207 FALLING_COUNTER.D.13 DC 0
V363 FALLING_COMP.Q_b FALLING_COMP.INV_Q.O DC 0
V364 FALLING_COMP.INV_Q.I FALLING_COMP.Q DC 0
V365 RISING_COUNTER.D.14 87 DC 0
V366 208 RISING_COUNTER.O.14 DC 0
V367 RISING_COUNTER.RSTb RISING_COUNTER.RST_INV.O DC 0
V368 RISING_COUNTER.RST_INV.I RISING_COUNTER.RST DC 0
V369 RISING_COUNTER.O.0 RISING_COUNTER.COUNT_DFF.Q DC 0
V370 RISING_COUNTER.COUNT_DFF.RSTb RISING_COUNTER.RSTb DC 0
V371 RISING_COUNTER.COUNT_DFF.D RISING_COUNTER.D.0 DC 0
V372 RISING_COUNTER.COUNT_DFF.CLK RISING_COUNTER.CLK DC 0
V373 RISING_COUNTER.D.0 59 DC 0
V374 209 RISING_COUNTER.O.0 DC 0
V375 RISING_COUNTER.O.1 60 DC 0
V376 210 RISING_COUNTER.RSTb DC 0
V377 211 RISING_COUNTER.D.1 DC 0
V378 212 RISING_COUNTER.D.0 DC 0
V379 RISING_COUNTER.D.1 61 DC 0
V380 213 RISING_COUNTER.O.1 DC 0
V381 RISING_COUNTER.O.2 62 DC 0
V382 214 RISING_COUNTER.RSTb DC 0
V383 215 RISING_COUNTER.D.2 DC 0
V384 216 RISING_COUNTER.D.1 DC 0
V385 RISING_COUNTER.D.2 63 DC 0
V386 217 RISING_COUNTER.O.2 DC 0
V387 RISING_COUNTER.O.3 64 DC 0
V388 218 RISING_COUNTER.RSTb DC 0
V389 219 RISING_COUNTER.D.3 DC 0
V390 220 RISING_COUNTER.D.2 DC 0
V391 RISING_COUNTER.D.3 65 DC 0
V392 221 RISING_COUNTER.O.3 DC 0
V393 RISING_COUNTER.O.4 66 DC 0
V394 222 RISING_COUNTER.RSTb DC 0
V395 223 RISING_COUNTER.D.4 DC 0
V396 224 RISING_COUNTER.D.3 DC 0
V397 RISING_COUNTER.D.4 67 DC 0
V398 225 RISING_COUNTER.O.4 DC 0
V399 RISING_COUNTER.O.5 68 DC 0
V400 226 RISING_COUNTER.RSTb DC 0
V401 227 RISING_COUNTER.D.5 DC 0
V402 228 RISING_COUNTER.D.4 DC 0
V403 RISING_COUNTER.D.5 69 DC 0
V404 229 RISING_COUNTER.O.5 DC 0
V405 RISING_COUNTER.O.6 70 DC 0
V406 230 RISING_COUNTER.RSTb DC 0
V407 231 RISING_COUNTER.D.6 DC 0
V408 232 RISING_COUNTER.D.5 DC 0
V409 RISING_COUNTER.D.6 71 DC 0
V410 233 RISING_COUNTER.O.6 DC 0
V411 RISING_COUNTER.O.7 72 DC 0
V412 234 RISING_COUNTER.RSTb DC 0
V413 235 RISING_COUNTER.D.7 DC 0
V414 236 RISING_COUNTER.D.6 DC 0
V415 RISING_COUNTER.D.7 73 DC 0
V416 237 RISING_COUNTER.O.7 DC 0
V417 RISING_COUNTER.O.8 74 DC 0
V418 238 RISING_COUNTER.RSTb DC 0
V419 239 RISING_COUNTER.D.8 DC 0
V420 240 RISING_COUNTER.D.7 DC 0
V421 RISING_COUNTER.D.8 75 DC 0
V422 241 RISING_COUNTER.O.8 DC 0
V423 RISING_COUNTER.O.9 76 DC 0
V424 242 RISING_COUNTER.RSTb DC 0
V425 243 RISING_COUNTER.D.9 DC 0
V426 244 RISING_COUNTER.D.8 DC 0
V427 RISING_COUNTER.D.9 77 DC 0
V428 245 RISING_COUNTER.O.9 DC 0
V429 RISING_COUNTER.O.10 78 DC 0
V430 246 RISING_COUNTER.RSTb DC 0
V431 247 RISING_COUNTER.D.10 DC 0
V432 248 RISING_COUNTER.D.9 DC 0
V433 RISING_COUNTER.D.10 79 DC 0
V434 249 RISING_COUNTER.O.10 DC 0
V435 RISING_COUNTER.O.11 80 DC 0
V436 250 RISING_COUNTER.RSTb DC 0
V437 251 RISING_COUNTER.D.11 DC 0
V438 252 RISING_COUNTER.D.10 DC 0
V439 RISING_COUNTER.D.11 81 DC 0
V440 253 RISING_COUNTER.O.11 DC 0
V441 RISING_COUNTER.O.12 82 DC 0
V442 254 RISING_COUNTER.RSTb DC 0
V443 255 RISING_COUNTER.D.12 DC 0
V444 256 RISING_COUNTER.D.11 DC 0
V445 RISING_COUNTER.D.12 83 DC 0
V446 257 RISING_COUNTER.O.12 DC 0
V447 RISING_COUNTER.O.13 84 DC 0
V448 258 RISING_COUNTER.RSTb DC 0
V449 259 RISING_COUNTER.D.13 DC 0
V450 260 RISING_COUNTER.D.12 DC 0
V451 RISING_COUNTER.D.13 85 DC 0
V452 261 RISING_COUNTER.O.13 DC 0
V453 RISING_COUNTER.O.14 86 DC 0
V454 262 RISING_COUNTER.RSTb DC 0
V455 263 RISING_COUNTER.D.14 DC 0
V456 264 RISING_COUNTER.D.13 DC 0
V457 FALLING_COUNTER.D.15 135 DC 0
V458 265 FALLING_COUNTER.O.15 DC 0
V459 FALLING_COUNTER.O.15 134 DC 0
V460 266 FALLING_COUNTER.RSTb DC 0
V461 267 FALLING_COUNTER.D.15 DC 0
V462 268 FALLING_COUNTER.D.14 DC 0
V463 FULL_COUNTER.D.18 37 DC 0
V464 269 FULL_COUNTER.O.18 DC 0
V465 FULL_COUNTER.RSTb FULL_COUNTER.RST_INV.O DC 0
V466 FULL_COUNTER.RST_INV.I FULL_COUNTER.RST DC 0
V467 FULL_COUNTER.O.0 FULL_COUNTER.COUNT_DFF.Q DC 0
V468 FULL_COUNTER.COUNT_DFF.RSTb FULL_COUNTER.RSTb DC 0
V469 FULL_COUNTER.COUNT_DFF.D FULL_COUNTER.D.0 DC 0
V470 FULL_COUNTER.COUNT_DFF.CLK FULL_COUNTER.CLK DC 0
V471 FULL_COUNTER.D.0 1 DC 0
V472 270 FULL_COUNTER.O.0 DC 0
V473 FULL_COUNTER.O.1 2 DC 0
V474 271 FULL_COUNTER.RSTb DC 0
V475 272 FULL_COUNTER.D.1 DC 0
V476 273 FULL_COUNTER.D.0 DC 0
V477 FULL_COUNTER.D.1 3 DC 0
V478 274 FULL_COUNTER.O.1 DC 0
V479 FULL_COUNTER.O.2 4 DC 0
V480 275 FULL_COUNTER.RSTb DC 0
V481 276 FULL_COUNTER.D.2 DC 0
V482 277 FULL_COUNTER.D.1 DC 0
V483 FULL_COUNTER.D.2 5 DC 0
V484 278 FULL_COUNTER.O.2 DC 0
V485 FULL_COUNTER.O.3 6 DC 0
V486 279 FULL_COUNTER.RSTb DC 0
V487 280 FULL_COUNTER.D.3 DC 0
V488 281 FULL_COUNTER.D.2 DC 0
V489 FULL_COUNTER.D.3 7 DC 0
V490 282 FULL_COUNTER.O.3 DC 0
V491 FULL_COUNTER.O.4 8 DC 0
V492 283 FULL_COUNTER.RSTb DC 0
V493 284 FULL_COUNTER.D.4 DC 0
V494 285 FULL_COUNTER.D.3 DC 0
V495 FULL_COUNTER.D.4 9 DC 0
V496 286 FULL_COUNTER.O.4 DC 0
V497 FULL_COUNTER.O.5 10 DC 0
V498 287 FULL_COUNTER.RSTb DC 0
V499 288 FULL_COUNTER.D.5 DC 0
V500 289 FULL_COUNTER.D.4 DC 0
V501 FULL_COUNTER.D.5 11 DC 0
V502 290 FULL_COUNTER.O.5 DC 0
V503 FULL_COUNTER.O.6 12 DC 0
V504 291 FULL_COUNTER.RSTb DC 0
V505 292 FULL_COUNTER.D.6 DC 0
V506 293 FULL_COUNTER.D.5 DC 0
V507 FULL_COUNTER.D.6 13 DC 0
V508 294 FULL_COUNTER.O.6 DC 0
V509 FULL_COUNTER.O.7 14 DC 0
V510 295 FULL_COUNTER.RSTb DC 0
V511 296 FULL_COUNTER.D.7 DC 0
V512 297 FULL_COUNTER.D.6 DC 0
V513 FULL_COUNTER.D.7 15 DC 0
V514 298 FULL_COUNTER.O.7 DC 0
V515 FULL_COUNTER.O.8 16 DC 0
V516 299 FULL_COUNTER.RSTb DC 0
V517 300 FULL_COUNTER.D.8 DC 0
V518 301 FULL_COUNTER.D.7 DC 0
V519 FULL_COUNTER.D.8 17 DC 0
V520 302 FULL_COUNTER.O.8 DC 0
V521 FULL_COUNTER.O.9 18 DC 0
V522 303 FULL_COUNTER.RSTb DC 0
V523 304 FULL_COUNTER.D.9 DC 0
V524 305 FULL_COUNTER.D.8 DC 0
V525 FULL_COUNTER.D.9 19 DC 0
V526 306 FULL_COUNTER.O.9 DC 0
V527 FULL_COUNTER.O.10 20 DC 0
V528 307 FULL_COUNTER.RSTb DC 0
V529 308 FULL_COUNTER.D.10 DC 0
V530 309 FULL_COUNTER.D.9 DC 0
V531 FULL_COUNTER.D.10 21 DC 0
V532 310 FULL_COUNTER.O.10 DC 0
V533 FULL_COUNTER.O.11 22 DC 0
V534 311 FULL_COUNTER.RSTb DC 0
V535 312 FULL_COUNTER.D.11 DC 0
V536 313 FULL_COUNTER.D.10 DC 0
V537 FULL_COUNTER.D.11 23 DC 0
V538 314 FULL_COUNTER.O.11 DC 0
V539 FULL_COUNTER.O.12 24 DC 0
V540 315 FULL_COUNTER.RSTb DC 0
V541 316 FULL_COUNTER.D.12 DC 0
V542 317 FULL_COUNTER.D.11 DC 0
V543 FULL_COUNTER.D.12 25 DC 0
V544 318 FULL_COUNTER.O.12 DC 0
V545 FULL_COUNTER.O.13 26 DC 0
V546 319 FULL_COUNTER.RSTb DC 0
V547 320 FULL_COUNTER.D.13 DC 0
V548 321 FULL_COUNTER.D.12 DC 0
V549 FULL_COUNTER.D.13 27 DC 0
V550 322 FULL_COUNTER.O.13 DC 0
V551 FULL_COUNTER.O.14 28 DC 0
V552 323 FULL_COUNTER.RSTb DC 0
V553 324 FULL_COUNTER.D.14 DC 0
V554 325 FULL_COUNTER.D.13 DC 0
V555 FULL_COUNTER.D.14 29 DC 0
V556 326 FULL_COUNTER.O.14 DC 0
V557 FULL_COUNTER.O.15 30 DC 0
V558 327 FULL_COUNTER.RSTb DC 0
V559 328 FULL_COUNTER.D.15 DC 0
V560 329 FULL_COUNTER.D.14 DC 0
V561 FULL_COUNTER.D.15 31 DC 0
V562 330 FULL_COUNTER.O.15 DC 0
V563 FULL_COUNTER.O.16 32 DC 0
V564 331 FULL_COUNTER.RSTb DC 0
V565 332 FULL_COUNTER.D.16 DC 0
V566 333 FULL_COUNTER.D.15 DC 0
V567 FULL_COUNTER.D.16 33 DC 0
V568 334 FULL_COUNTER.O.16 DC 0
V569 FULL_COUNTER.O.17 34 DC 0
V570 335 FULL_COUNTER.RSTb DC 0
V571 336 FULL_COUNTER.D.17 DC 0
V572 337 FULL_COUNTER.D.16 DC 0
V573 FULL_COUNTER.D.17 35 DC 0
V574 338 FULL_COUNTER.O.17 DC 0
V575 FULL_COUNTER.O.18 36 DC 0
V576 339 FULL_COUNTER.RSTb DC 0
V577 340 FULL_COUNTER.D.18 DC 0
V578 341 FULL_COUNTER.D.17 DC 0
V579 RISING_COUNTER.D.15 89 DC 0
V580 342 RISING_COUNTER.O.15 DC 0
V581 RISING_COUNTER.O.15 88 DC 0
V582 343 RISING_COUNTER.RSTb DC 0
V583 344 RISING_COUNTER.D.15 DC 0
V584 345 RISING_COUNTER.D.14 DC 0
V585 FULL_COUNTER.D.19 39 DC 0
V586 346 FULL_COUNTER.O.19 DC 0
V587 FULL_COUNTER.O.19 38 DC 0
V588 347 FULL_COUNTER.RSTb DC 0
V589 348 FULL_COUNTER.D.19 DC 0
V590 349 FULL_COUNTER.D.18 DC 0
V591 CLOCK_GEN.SR_OE.Qb CLOCK_GEN.SR_OE.NANDQb.O DC 0
V592 CLOCK_GEN.SR_OE.NANDQb.B CLOCK_GEN.SR_OE.Q DC 0
V593 CLOCK_GEN.SR_OE.NANDQb.A CLOCK_GEN.SR_OE.Rb DC 0
V594 CLOCK_GEN.SR_OE.Q CLOCK_GEN.SR_OE.NANDQ.O DC 0
V595 CLOCK_GEN.SR_OE.NANDQ.B CLOCK_GEN.SR_OE.Qb DC 0
V596 CLOCK_GEN.SR_OE.NANDQ.A CLOCK_GEN.SR_OE.Sb DC 0
V597 FALLING_COMP.SR_MEM.Q FALLING_COMP.SR_MEM.NANDQ.O DC 0
V598 FALLING_COMP.SR_MEM.NANDQ.B FALLING_COMP.SR_MEM.Qb DC 0
V599 FALLING_COMP.SR_MEM.NANDQ.A FALLING_COMP.SR_MEM.Sb DC 0
V600 FALLING_COMP.SR_MEM.Qb FALLING_COMP.SR_MEM.NANDQb.O DC 0
V601 FALLING_COMP.SR_MEM.NANDQb.B FALLING_COMP.SR_MEM.Q DC 0
V602 FALLING_COMP.SR_MEM.NANDQb.A FALLING_COMP.SR_MEM.Rb DC 0
V603 FINISH_COMP.SR_MEM.Q FINISH_COMP.SR_MEM.NANDQ.O DC 0
V604 FINISH_COMP.SR_MEM.NANDQ.B FINISH_COMP.SR_MEM.Qb DC 0
V605 FINISH_COMP.SR_MEM.NANDQ.A FINISH_COMP.SR_MEM.Sb DC 0
V606 FINISH_COMP.SR_MEM.Qb FINISH_COMP.SR_MEM.NANDQb.O DC 0
V607 FINISH_COMP.SR_MEM.NANDQb.B FINISH_COMP.SR_MEM.Q DC 0
V608 FINISH_COMP.SR_MEM.NANDQb.A FINISH_COMP.SR_MEM.Rb DC 0
V609 CLOCK_GEN.SR_Op.Qb CLOCK_GEN.SR_Op.NANDQb.O DC 0
V610 CLOCK_GEN.SR_Op.NANDQb.B CLOCK_GEN.SR_Op.Q DC 0
V611 CLOCK_GEN.SR_Op.NANDQb.A CLOCK_GEN.SR_Op.Rb DC 0
V612 CLOCK_GEN.SR_Op.Q CLOCK_GEN.SR_Op.NANDQ.O DC 0
V613 CLOCK_GEN.SR_Op.NANDQ.B CLOCK_GEN.SR_Op.Qb DC 0
V614 CLOCK_GEN.SR_Op.NANDQ.A CLOCK_GEN.SR_Op.Sb DC 0
V615 RISING_COMP.SR_MEM.Q RISING_COMP.SR_MEM.NANDQ.O DC 0
V616 RISING_COMP.SR_MEM.NANDQ.B RISING_COMP.SR_MEM.Qb DC 0
V617 RISING_COMP.SR_MEM.NANDQ.A RISING_COMP.SR_MEM.Sb DC 0
V618 RISING_COMP.SR_MEM.Qb RISING_COMP.SR_MEM.NANDQb.O DC 0
V619 RISING_COMP.SR_MEM.NANDQb.B RISING_COMP.SR_MEM.Q DC 0
V620 RISING_COMP.SR_MEM.NANDQb.A RISING_COMP.SR_MEM.Rb DC 0
.ends