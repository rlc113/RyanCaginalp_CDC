`include "Physical_Gates.v"

`ifndef INVCHAIN_GUARD
`define INVCHAIN_GUARD

module Normal_Inverter_Chain(input I, output O);
endmodule


module Cap_Inverter_Chain(input I, output O);
endmodule


module Finish_Inverter_Chain(input I, output Ob, output O);
endmodule

`endif