`include "Physical_Gates.v"

`ifndef CHAIN_DRIVER_GUARD
`define CHAIN_DRIVER_GUARD

module chain_driver(input Next_Edge_LowV, output Next_Edge_HighV);
endmodule

`endif