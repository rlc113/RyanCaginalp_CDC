.subckt CDC Reset Next_Edge_HighV Falling_Y Rising_Y Conversion_Finished V_GND V_LOW V_HIGH V_SENSE Falling_Low Falling_Cap Finish_Delay FALLING_COMP.Qb_b FALLING_COMP.Db_Plus FALLING_COMP.Output_Enable FALLING_COMP.Y


X0 CLOCK_GEN.INV_R.O CLOCK_GEN.SR_Op.Q CLOCK_GEN.SR_Op.Qb sky130_fd_sc_hd__nand2_8
X1 FINISH_COMP.INV_DM.O FINISH_COMP.SR_MEM.Q FINISH_COMP.SR_MEM.Qb sky130_fd_sc_hd__nand2_8
X2 RISING_COMP.INV_DM.O RISING_COMP.SR_MEM.Q RISING_COMP.SR_MEM.Qb sky130_fd_sc_hd__nand2_8
X3 CLOCK_GEN.NAND_DR.O CLOCK_GEN.SR_OE.Q CLOCK_GEN.SR_OE.Qb sky130_fd_sc_hd__nand2_8
X4 FALLING_COMP.INV_DM.O FALLING_COMP.SR_MEM.Q FALLING_COMP.SR_MEM.Qb sky130_fd_sc_hd__nand2_8
X5 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_INV0.O sky130_fd_sc_hd__inv_1
X6 FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_INV1.O sky130_fd_sc_hd__inv_1
X7 FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_INV2.O sky130_fd_sc_hd__inv_1
X8 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_INV3.O sky130_fd_sc_hd__inv_1
X9 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_INV4.O sky130_fd_sc_hd__inv_1
X10 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_INV5.O sky130_fd_sc_hd__inv_1
X11 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_INV6.O sky130_fd_sc_hd__inv_1
X12 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_INV7.O sky130_fd_sc_hd__inv_1
X13 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_INV8.O sky130_fd_sc_hd__inv_1
X14 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_INV9.O sky130_fd_sc_hd__inv_1
X15 FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_INV10.O sky130_fd_sc_hd__inv_1
X16 FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_INV11.O sky130_fd_sc_hd__inv_1
X17 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_INV12.O sky130_fd_sc_hd__inv_1
X18 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_INV13.O sky130_fd_sc_hd__inv_1
X19 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_INV14.O sky130_fd_sc_hd__inv_1
X20 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_INV15.O sky130_fd_sc_hd__inv_1
X21 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_INV16.O sky130_fd_sc_hd__inv_1
X22 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_INV17.O sky130_fd_sc_hd__inv_1
X23 FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_INV18.O sky130_fd_sc_hd__inv_1
X24 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_INV19.O sky130_fd_sc_hd__inv_1
X25 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_INV0.O CLOCK_GEN.NOT_CLK.O FULL_COUNTER.COUNT_SUB_DFF0.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X26 FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_INV1.O FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF1.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X27 FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_INV2.O FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF2.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X28 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_INV3.O FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF3.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X29 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_INV4.O FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF4.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X30 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_INV5.O FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF5.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X31 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_INV6.O FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF6.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X32 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_INV7.O FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF7.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X33 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_INV8.O FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF8.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X34 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_INV9.O FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF9.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X35 FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_INV10.O FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF10.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X36 FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_INV11.O FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_DFF11.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X37 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_INV12.O FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_DFF12.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X38 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_INV13.O FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF13.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X39 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_INV14.O FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF14.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X40 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_INV15.O FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF15.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X41 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_INV16.O FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF16.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X42 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_INV17.O FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF17.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X43 FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_INV18.O FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF18.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X44 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_INV19.O FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_DFF19.Qb FULL_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X45 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_INV0.O sky130_fd_sc_hd__inv_1
X46 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_INV1.O sky130_fd_sc_hd__inv_1
X47 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_INV2.O sky130_fd_sc_hd__inv_1
X48 RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_INV3.O sky130_fd_sc_hd__inv_1
X49 RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_INV4.O sky130_fd_sc_hd__inv_1
X50 RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_INV5.O sky130_fd_sc_hd__inv_1
X51 RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_INV6.O sky130_fd_sc_hd__inv_1
X52 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_INV7.O sky130_fd_sc_hd__inv_1
X53 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_INV8.O sky130_fd_sc_hd__inv_1
X54 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_INV9.O sky130_fd_sc_hd__inv_1
X55 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_INV10.O sky130_fd_sc_hd__inv_1
X56 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_INV11.O sky130_fd_sc_hd__inv_1
X57 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_INV12.O sky130_fd_sc_hd__inv_1
X58 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_INV13.O sky130_fd_sc_hd__inv_1
X59 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_INV14.O sky130_fd_sc_hd__inv_1
X60 RISING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_INV15.O sky130_fd_sc_hd__inv_1
X61 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_INV0.O RISING_COMP.NAND3_COMP.O RISING_COUNTER.COUNT_SUB_DFF0.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X62 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_INV1.O RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF1.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X63 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_INV2.O RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF2.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X64 RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_INV3.O RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF3.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X65 RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_INV4.O RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF4.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X66 RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_INV5.O RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF5.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X67 RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_INV6.O RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF6.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X68 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_INV7.O RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF7.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X69 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_INV8.O RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF8.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X70 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_INV9.O RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF9.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X71 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_INV10.O RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF10.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X72 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_INV11.O RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF11.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X73 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_INV12.O RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF12.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X74 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_INV13.O RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF13.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X75 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_INV14.O RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF14.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X76 RISING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_INV15.O RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF15.Qb RISING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X77 FALLING_COUNTER.COUNT_SUB_DFF0.Q FALLING_COUNTER.COUNT_SUB_INV0.O sky130_fd_sc_hd__inv_1
X78 FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_INV1.O sky130_fd_sc_hd__inv_1
X79 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_INV2.O sky130_fd_sc_hd__inv_1
X80 FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_INV3.O sky130_fd_sc_hd__inv_1
X81 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_INV4.O sky130_fd_sc_hd__inv_1
X82 FALLING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_INV5.O sky130_fd_sc_hd__inv_1
X83 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_INV6.O sky130_fd_sc_hd__inv_1
X84 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_INV7.O sky130_fd_sc_hd__inv_1
X85 FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_INV8.O sky130_fd_sc_hd__inv_1
X86 FALLING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_INV9.O sky130_fd_sc_hd__inv_1
X87 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_INV10.O sky130_fd_sc_hd__inv_1
X88 FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_INV11.O sky130_fd_sc_hd__inv_1
X89 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_INV12.O sky130_fd_sc_hd__inv_1
X90 FALLING_COUNTER.COUNT_SUB_DFF13.Q FALLING_COUNTER.COUNT_SUB_INV13.O sky130_fd_sc_hd__inv_1
X91 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_INV14.O sky130_fd_sc_hd__inv_1
X92 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_INV15.O sky130_fd_sc_hd__inv_1
X93 FALLING_COUNTER.COUNT_SUB_DFF0.Q FALLING_COUNTER.COUNT_SUB_INV0.O FALLING_COMP.NAND3_COMP.O FALLING_COUNTER.COUNT_SUB_DFF0.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X94 FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_INV1.O FALLING_COUNTER.COUNT_SUB_DFF0.Q FALLING_COUNTER.COUNT_SUB_DFF1.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X95 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_INV2.O FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_DFF2.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X96 FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_INV3.O FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF3.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X97 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_INV4.O FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_DFF4.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X98 FALLING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_INV5.O FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF5.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X99 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_INV6.O FALLING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_DFF6.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X100 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_INV7.O FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF7.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X101 FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_INV8.O FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF8.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X102 FALLING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_INV9.O FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF9.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X103 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_INV10.O FALLING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF10.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X104 FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_INV11.O FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF11.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X105 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_INV12.O FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF12.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X106 FALLING_COUNTER.COUNT_SUB_DFF13.Q FALLING_COUNTER.COUNT_SUB_INV13.O FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF13.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X107 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_INV14.O FALLING_COUNTER.COUNT_SUB_DFF13.Q FALLING_COUNTER.COUNT_SUB_DFF14.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X108 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_INV15.O FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF15.Qb FALLING_COUNTER.RSTb V_LOW sky130_fd_sc_hd__dfbbn_1
X109 LOW_CHAIN.low_chain_inv1.O LOW_CHAIN.low_chain_inv2.O sky130_fd_sc_hd__inv_1
X110 LOW_CHAIN.low_chain_inv2.O LOW_CHAIN.low_chain_inv3.O sky130_fd_sc_hd__inv_1
X111 LOW_CHAIN.low_chain_inv3.O LOW_CHAIN.low_chain_inv4.O sky130_fd_sc_hd__inv_1
X112 LOW_CHAIN.low_chain_inv4.O LOW_CHAIN.low_chain_inv5.O sky130_fd_sc_hd__inv_1
X113 LOW_CHAIN.low_chain_inv5.O LOW_CHAIN.low_chain_inv6.O sky130_fd_sc_hd__inv_1
X114 LOW_CHAIN.low_chain_inv6.O LOW_CHAIN.low_chain_inv7.O sky130_fd_sc_hd__inv_1
X115 LOW_CHAIN.low_chain_inv7.O LOW_CHAIN.low_chain_inv8.O sky130_fd_sc_hd__inv_1
X116 LOW_CHAIN.low_chain_inv8.O LOW_CHAIN.low_chain_inv9.O sky130_fd_sc_hd__inv_1
X117 LOW_CHAIN.low_chain_inv9.O LOW_CHAIN.low_chain_inv10.O sky130_fd_sc_hd__inv_1
X118 LOW_CHAIN.low_chain_inv10.O LOW_CHAIN.low_chain_inv11.O sky130_fd_sc_hd__inv_1
X119 LOW_CHAIN.low_chain_inv11.O LOW_CHAIN.low_chain_inv12.O sky130_fd_sc_hd__inv_1
X120 LOW_CHAIN.low_chain_inv12.O LOW_CHAIN.low_chain_inv13.O sky130_fd_sc_hd__inv_1
X121 LOW_CHAIN.low_chain_inv13.O LOW_CHAIN.low_chain_inv14.O sky130_fd_sc_hd__inv_1
X122 LOW_CHAIN.low_chain_inv14.O LOW_CHAIN.low_chain_inv15.O sky130_fd_sc_hd__inv_1
X123 LOW_CHAIN.low_chain_inv15.O LOW_CHAIN.low_chain_inv16.O sky130_fd_sc_hd__inv_1
X124 FINISH_CHAIN.finish_chain_inv15.O CLOCK_GEN.INV_F.O sky130_fd_sc_hd__inv_1
X125 FALLING_COMP.NAND2_COMP.O CLOCK_GEN.INV_F.O CLOCK_GEN.NAND_DF.O sky130_fd_sc_hd__nand2_1
X126 CLOCK_GEN.NAND_DF.O CLOCK_GEN.SR_OE.Qb CLOCK_GEN.SR_OE.Q sky130_fd_sc_hd__nand2_8
X127 CLOCK_GEN.SR_OE.Q CLOCK_GEN.INV_OE.O sky130_fd_sc_hd__inv_1
X128 Reset CLOCK_GEN.INV_R.O sky130_fd_sc_hd__inv_1
X129 FINISH_COMP.NAND3_COMP.O CLOCK_GEN.SR_Op.Qb CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand2_8
X130 Reset CLOCK_GEN.SR_Op.Q CLOCK_GEN.NOR_CLK.O sky130_fd_sc_hd__nor2_1
X131 CLOCK_GEN.SR_OE.Q CLOCK_GEN.NOR_CLK.O CLOCK_GEN.NAND_CLK.O sky130_fd_sc_hd__nand2_1
X132 CLOCK_GEN.NAND_CLK.O CLOCK_GEN.NOT_CLK.O sky130_fd_sc_hd__inv_1
X133 FINISH_CHAIN.finish_chain_inv16.O FINISH_COMP.INV_DM.O sky130_fd_sc_hd__inv_1
X134 FINISH_COMP.INV_DP.O FINISH_COMP.SR_MEM.Qb FINISH_COMP.SR_MEM.Q sky130_fd_sc_hd__nand2_8
X135 FINISH_COMP.SR_MEM.Q FINISH_COMP.INV_Q.O sky130_fd_sc_hd__inv_1
X136 FINISH_COMP.SR_MEM.Qb FINISH_COMP.INV_Qb.O sky130_fd_sc_hd__inv_1
X137 INV_RISING_CAP.O FINISH_CHAIN.finish_chain_inv16.O FINISH_COMP.NAND2_COMP.O sky130_fd_sc_hd__nand2_1
X138 FINISH_COMP.INV_Qb.O FINISH_COMP.INV_DP.O FINISH_COMP.NAND3_COMP.O CLOCK_GEN.INV_OE.O sky130_fd_sc_hd__nand3_1
X139 INV_RISING_LOW.O RISING_COMP.INV_DM.O sky130_fd_sc_hd__inv_1
X140 RISING_COMP.INV_DP.O RISING_COMP.SR_MEM.Qb RISING_COMP.SR_MEM.Q sky130_fd_sc_hd__nand2_8
X141 RISING_COMP.SR_MEM.Q RISING_COMP.INV_Q.O sky130_fd_sc_hd__inv_1
X142 RISING_COMP.SR_MEM.Qb RISING_COMP.INV_Qb.O sky130_fd_sc_hd__inv_1
X143 INV_RISING_CAP.O INV_RISING_LOW.O RISING_COMP.NAND2_COMP.O sky130_fd_sc_hd__nand2_1
X144 RISING_COMP.INV_Qb.O RISING_COMP.INV_DP.O RISING_COMP.NAND3_COMP.O CLOCK_GEN.INV_OE.O sky130_fd_sc_hd__nand3_1
X145 LOW_CHAIN.low_chain_inv16.O FALLING_COMP.INV_DM.O sky130_fd_sc_hd__inv_1
X146 FALLING_COMP.INV_DP.O FALLING_COMP.SR_MEM.Qb FALLING_COMP.SR_MEM.Q sky130_fd_sc_hd__nand2_8
X147 FALLING_COMP.SR_MEM.Q FALLING_COMP.INV_Q.O sky130_fd_sc_hd__inv_1
X148 FALLING_COMP.SR_MEM.Qb FALLING_COMP.INV_Qb.O sky130_fd_sc_hd__inv_1
X149 CAP_CHAIN.cap_chain_inv16.O LOW_CHAIN.low_chain_inv16.O FALLING_COMP.NAND2_COMP.O sky130_fd_sc_hd__nand2_1
X150 FALLING_COMP.INV_Qb.O FALLING_COMP.INV_DP.O FALLING_COMP.NAND3_COMP.O CLOCK_GEN.SR_OE.Q sky130_fd_sc_hd__nand3_1
X151 CAP_CHAIN.cap_chain_inv1.O CAP_CHAIN.cap_chain_inv2.O sky130_fd_sc_hd__inv_1
X152 CAP_CHAIN.cap_chain_inv2.O CAP_CHAIN.cap_chain_inv3.O sky130_fd_sc_hd__inv_1
X153 CAP_CHAIN.cap_chain_inv3.O CAP_CHAIN.cap_chain_inv4.O sky130_fd_sc_hd__inv_1
X154 CAP_CHAIN.cap_chain_inv4.O CAP_CHAIN.cap_chain_inv5.O sky130_fd_sc_hd__inv_1
X155 CAP_CHAIN.cap_chain_inv5.O CAP_CHAIN.cap_chain_inv6.O sky130_fd_sc_hd__inv_1
X156 CAP_CHAIN.cap_chain_inv6.O CAP_CHAIN.cap_chain_inv7.O sky130_fd_sc_hd__inv_1
X157 CAP_CHAIN.cap_chain_inv7.O CAP_CHAIN.cap_chain_inv8.O sky130_fd_sc_hd__inv_1
X158 CAP_CHAIN.cap_chain_inv8.O CAP_CHAIN.cap_chain_inv9.O sky130_fd_sc_hd__inv_1
X159 CAP_CHAIN.cap_chain_inv9.O CAP_CHAIN.cap_chain_inv10.O sky130_fd_sc_hd__inv_1
X160 CAP_CHAIN.cap_chain_inv10.O CAP_CHAIN.cap_chain_inv11.O sky130_fd_sc_hd__inv_1
X161 CAP_CHAIN.cap_chain_inv11.O CAP_CHAIN.cap_chain_inv12.O sky130_fd_sc_hd__inv_1
X162 CAP_CHAIN.cap_chain_inv12.O CAP_CHAIN.cap_chain_inv13.O sky130_fd_sc_hd__inv_1
X163 CAP_CHAIN.cap_chain_inv13.O CAP_CHAIN.cap_chain_inv14.O sky130_fd_sc_hd__inv_1
X164 CAP_CHAIN.cap_chain_inv14.O CAP_CHAIN.cap_chain_inv15.O sky130_fd_sc_hd__inv_1
X165 CAP_CHAIN.cap_chain_inv15.O CAP_CHAIN.cap_chain_inv16.O sky130_fd_sc_hd__inv_1
X166 FINISH_CHAIN.finish_chain_inv1.O FINISH_CHAIN.finish_chain_inv2.O sky130_fd_sc_hd__inv_1
X167 FINISH_CHAIN.finish_chain_inv2.O FINISH_CHAIN.finish_chain_inv3.O sky130_fd_sc_hd__inv_1
X168 FINISH_CHAIN.finish_chain_inv3.O FINISH_CHAIN.finish_chain_inv4.O sky130_fd_sc_hd__inv_1
X169 FINISH_CHAIN.finish_chain_inv4.O FINISH_CHAIN.finish_chain_inv5.O sky130_fd_sc_hd__inv_1
X170 FINISH_CHAIN.finish_chain_inv5.O FINISH_CHAIN.finish_chain_inv6.O sky130_fd_sc_hd__inv_1
X171 FINISH_CHAIN.finish_chain_inv6.O FINISH_CHAIN.finish_chain_inv7.O sky130_fd_sc_hd__inv_1
X172 FINISH_CHAIN.finish_chain_inv7.O FINISH_CHAIN.finish_chain_inv8.O sky130_fd_sc_hd__inv_1
X173 FINISH_CHAIN.finish_chain_inv8.O FINISH_CHAIN.finish_chain_inv9.O sky130_fd_sc_hd__inv_1
X174 FINISH_CHAIN.finish_chain_inv9.O FINISH_CHAIN.finish_chain_inv10.O sky130_fd_sc_hd__inv_1
X175 FINISH_CHAIN.finish_chain_inv10.O FINISH_CHAIN.finish_chain_inv11.O sky130_fd_sc_hd__inv_1
X176 FINISH_CHAIN.finish_chain_inv11.O FINISH_CHAIN.finish_chain_inv12.O sky130_fd_sc_hd__inv_1
X177 FINISH_CHAIN.finish_chain_inv12.O FINISH_CHAIN.finish_chain_inv13.O sky130_fd_sc_hd__inv_1
X178 FINISH_CHAIN.finish_chain_inv13.O FINISH_CHAIN.finish_chain_inv14.O sky130_fd_sc_hd__inv_1
X179 FINISH_CHAIN.finish_chain_inv14.O FINISH_CHAIN.finish_chain_inv15.O sky130_fd_sc_hd__inv_1
X180 FINISH_CHAIN.finish_chain_inv15.O FINISH_CHAIN.finish_chain_inv16.O sky130_fd_sc_hd__inv_1
X181 V_HIGH Reset V_SENSE transmission_gate
X182 Next_Edge_LowV_b Next_Edge_HighV sky130_fd_sc_hd__inv_2
X183 CLOCK_GEN.NOT_CLK.O Next_Edge_LowV_b sky130_fd_sc_hd__inv_1
X184 Reset FULL_COUNTER.RSTb sky130_fd_sc_hd__inv_16
X185 RISING_COMP.NAND2_COMP.O FINISH_CHAIN.finish_chain_inv15.O CLOCK_GEN.NAND_DR.O sky130_fd_sc_hd__nand2_1
X186 INV_RISING_CAP.O FINISH_COMP.INV_DP.O sky130_fd_sc_hd__inv_1
X187 Reset RISING_COUNTER.RSTb sky130_fd_sc_hd__inv_16
X188 INV_RISING_CAP.O RISING_COMP.INV_DP.O sky130_fd_sc_hd__inv_1
X189 Reset FALLING_COUNTER.RSTb sky130_fd_sc_hd__inv_16
X190 CAP_CHAIN.cap_chain_inv16.O FALLING_COMP.INV_DP.O sky130_fd_sc_hd__inv_1
X191 INV_RISING_LOW.O FINISH_CHAIN.finish_chain_inv1.O sky130_fd_sc_hd__inv_1
X192 CAP_CHAIN.cap_chain_inv16.O INV_RISING_CAP.O sky130_fd_sc_hd__inv_1
X193 LOW_CHAIN.low_chain_inv16.O INV_RISING_LOW.O sky130_fd_sc_hd__inv_1
X194 Next_Edge_HighV CAP_CHAIN.cap_chain_inv1.O sky130_fd_sc_hd__inv_1
X195 Next_Edge_HighV LOW_CHAIN.low_chain_inv1.O sky130_fd_sc_hd__inv_1
V0 Rising_Low INV_RISING_LOW.O DC 0
V1 INV_RISING_LOW.I Falling_Low DC 0
V2 Finish_Low FINISH_CHAIN.O DC 0
V3 Finish_Delay FINISH_CHAIN.Ob DC 0
V4 FINISH_CHAIN.I Rising_Low DC 0
V5 Falling_Cap CAP_CHAIN.O DC 0
V6 CAP_CHAIN.I Next_Edge_HighV DC 0
V7 Falling_Y FALLING_COMP.Y DC 0
V8 Falling_Done FALLING_COMP.Done DC 0
V9 FALLING_COMP.Output_Enable Falling_Output_Enable DC 0
V10 FALLING_COMP.D_Minus Falling_Low DC 0
V11 FALLING_COMP.D_Plus Falling_Cap DC 0
V12 Rising_Cap INV_RISING_CAP.O DC 0
V13 INV_RISING_CAP.I Falling_Cap DC 0
V14 Rising_Y RISING_COMP.Y DC 0
V15 Rising_Done RISING_COMP.Done DC 0
V16 RISING_COMP.Output_Enable Rising_Output_Enable DC 0
V17 RISING_COMP.D_Minus Rising_Low DC 0
V18 RISING_COMP.D_Plus Rising_Cap DC 0
V19 Finish FINISH_COMP.Y DC 0
V20 FINISH_COMP.Output_Enable Rising_Output_Enable DC 0
V21 FINISH_COMP.D_Minus Finish_Low DC 0
V22 FINISH_COMP.D_Plus Rising_Cap DC 0
V23 Conversion_Finished CLOCK_GEN.Conv_Finish DC 0
V24 Next_Edge_LowV CLOCK_GEN.Next_Edge DC 0
V25 Falling_Output_Enable CLOCK_GEN.OE_Falling DC 0
V26 Rising_Output_Enable CLOCK_GEN.OE_Rising DC 0
V27 CLOCK_GEN.Finish Finish DC 0
V28 CLOCK_GEN.Reset Reset DC 0
V29 CLOCK_GEN.Finish_Delay Finish_Delay DC 0
V30 CLOCK_GEN.Done_Falling Falling_Done DC 0
V31 CLOCK_GEN.Done_Rising Rising_Done DC 0
V32 Falling_Low LOW_CHAIN.O DC 0
V33 LOW_CHAIN.I Next_Edge_HighV DC 0
V34 D_SUB2.0 FALLING_COUNTER.O.0 DC 0
V35 D_SUB2.1 FALLING_COUNTER.O.1 DC 0
V36 D_SUB2.2 FALLING_COUNTER.O.2 DC 0
V37 D_SUB2.3 FALLING_COUNTER.O.3 DC 0
V38 D_SUB2.4 FALLING_COUNTER.O.4 DC 0
V39 D_SUB2.5 FALLING_COUNTER.O.5 DC 0
V40 D_SUB2.6 FALLING_COUNTER.O.6 DC 0
V41 D_SUB2.7 FALLING_COUNTER.O.7 DC 0
V42 D_SUB2.8 FALLING_COUNTER.O.8 DC 0
V43 D_SUB2.9 FALLING_COUNTER.O.9 DC 0
V44 D_SUB2.10 FALLING_COUNTER.O.10 DC 0
V45 D_SUB2.11 FALLING_COUNTER.O.11 DC 0
V46 D_SUB2.12 FALLING_COUNTER.O.12 DC 0
V47 D_SUB2.13 FALLING_COUNTER.O.13 DC 0
V48 D_SUB2.14 FALLING_COUNTER.O.14 DC 0
V49 D_SUB2.15 FALLING_COUNTER.O.15 DC 0
V50 FALLING_COUNTER.RST Reset DC 0
V51 FALLING_COUNTER.CLK Falling_Y DC 0
V52 D_SUB1.0 RISING_COUNTER.O.0 DC 0
V53 D_SUB1.1 RISING_COUNTER.O.1 DC 0
V54 D_SUB1.2 RISING_COUNTER.O.2 DC 0
V55 D_SUB1.3 RISING_COUNTER.O.3 DC 0
V56 D_SUB1.4 RISING_COUNTER.O.4 DC 0
V57 D_SUB1.5 RISING_COUNTER.O.5 DC 0
V58 D_SUB1.6 RISING_COUNTER.O.6 DC 0
V59 D_SUB1.7 RISING_COUNTER.O.7 DC 0
V60 D_SUB1.8 RISING_COUNTER.O.8 DC 0
V61 D_SUB1.9 RISING_COUNTER.O.9 DC 0
V62 D_SUB1.10 RISING_COUNTER.O.10 DC 0
V63 D_SUB1.11 RISING_COUNTER.O.11 DC 0
V64 D_SUB1.12 RISING_COUNTER.O.12 DC 0
V65 D_SUB1.13 RISING_COUNTER.O.13 DC 0
V66 D_SUB1.14 RISING_COUNTER.O.14 DC 0
V67 D_SUB1.15 RISING_COUNTER.O.15 DC 0
V68 RISING_COUNTER.RST Reset DC 0
V69 RISING_COUNTER.CLK Rising_Y DC 0
V70 D_MAIN.0 FULL_COUNTER.O.0 DC 0
V71 D_MAIN.1 FULL_COUNTER.O.1 DC 0
V72 D_MAIN.2 FULL_COUNTER.O.2 DC 0
V73 D_MAIN.3 FULL_COUNTER.O.3 DC 0
V74 D_MAIN.4 FULL_COUNTER.O.4 DC 0
V75 D_MAIN.5 FULL_COUNTER.O.5 DC 0
V76 D_MAIN.6 FULL_COUNTER.O.6 DC 0
V77 D_MAIN.7 FULL_COUNTER.O.7 DC 0
V78 D_MAIN.8 FULL_COUNTER.O.8 DC 0
V79 D_MAIN.9 FULL_COUNTER.O.9 DC 0
V80 D_MAIN.10 FULL_COUNTER.O.10 DC 0
V81 D_MAIN.11 FULL_COUNTER.O.11 DC 0
V82 D_MAIN.12 FULL_COUNTER.O.12 DC 0
V83 D_MAIN.13 FULL_COUNTER.O.13 DC 0
V84 D_MAIN.14 FULL_COUNTER.O.14 DC 0
V85 D_MAIN.15 FULL_COUNTER.O.15 DC 0
V86 D_MAIN.16 FULL_COUNTER.O.16 DC 0
V87 D_MAIN.17 FULL_COUNTER.O.17 DC 0
V88 D_MAIN.18 FULL_COUNTER.O.18 DC 0
V89 D_MAIN.19 FULL_COUNTER.O.19 DC 0
V90 FULL_COUNTER.RST Reset DC 0
V91 FULL_COUNTER.CLK Next_Edge_LowV DC 0
V92 LOW_CHAIN.low_chain1 LOW_CHAIN.low_chain_inv1.O DC 0
V93 LOW_CHAIN.low_chain_inv1.I LOW_CHAIN.I DC 0
V94 LOW_CHAIN.low_chain2 LOW_CHAIN.low_chain_inv2.O DC 0
V95 LOW_CHAIN.low_chain_inv2.I LOW_CHAIN.low_chain1 DC 0
V96 LOW_CHAIN.low_chain3 LOW_CHAIN.low_chain_inv3.O DC 0
V97 LOW_CHAIN.low_chain_inv3.I LOW_CHAIN.low_chain2 DC 0
V98 LOW_CHAIN.low_chain4 LOW_CHAIN.low_chain_inv4.O DC 0
V99 LOW_CHAIN.low_chain_inv4.I LOW_CHAIN.low_chain3 DC 0
V100 LOW_CHAIN.low_chain5 LOW_CHAIN.low_chain_inv5.O DC 0
V101 LOW_CHAIN.low_chain_inv5.I LOW_CHAIN.low_chain4 DC 0
V102 LOW_CHAIN.low_chain6 LOW_CHAIN.low_chain_inv6.O DC 0
V103 LOW_CHAIN.low_chain_inv6.I LOW_CHAIN.low_chain5 DC 0
V104 LOW_CHAIN.low_chain7 LOW_CHAIN.low_chain_inv7.O DC 0
V105 LOW_CHAIN.low_chain_inv7.I LOW_CHAIN.low_chain6 DC 0
V106 LOW_CHAIN.low_chain8 LOW_CHAIN.low_chain_inv8.O DC 0
V107 LOW_CHAIN.low_chain_inv8.I LOW_CHAIN.low_chain7 DC 0
V108 LOW_CHAIN.low_chain9 LOW_CHAIN.low_chain_inv9.O DC 0
V109 LOW_CHAIN.low_chain_inv9.I LOW_CHAIN.low_chain8 DC 0
V110 LOW_CHAIN.low_chain10 LOW_CHAIN.low_chain_inv10.O DC 0
V111 LOW_CHAIN.low_chain_inv10.I LOW_CHAIN.low_chain9 DC 0
V112 LOW_CHAIN.low_chain11 LOW_CHAIN.low_chain_inv11.O DC 0
V113 LOW_CHAIN.low_chain_inv11.I LOW_CHAIN.low_chain10 DC 0
V114 LOW_CHAIN.low_chain12 LOW_CHAIN.low_chain_inv12.O DC 0
V115 LOW_CHAIN.low_chain_inv12.I LOW_CHAIN.low_chain11 DC 0
V116 LOW_CHAIN.low_chain13 LOW_CHAIN.low_chain_inv13.O DC 0
V117 LOW_CHAIN.low_chain_inv13.I LOW_CHAIN.low_chain12 DC 0
V118 LOW_CHAIN.low_chain14 LOW_CHAIN.low_chain_inv14.O DC 0
V119 LOW_CHAIN.low_chain_inv14.I LOW_CHAIN.low_chain13 DC 0
V120 LOW_CHAIN.low_chain15 LOW_CHAIN.low_chain_inv15.O DC 0
V121 LOW_CHAIN.low_chain_inv15.I LOW_CHAIN.low_chain14 DC 0
V122 LOW_CHAIN.O LOW_CHAIN.low_chain_inv16.O DC 0
V123 LOW_CHAIN.low_chain_inv16.I LOW_CHAIN.low_chain15 DC 0
V124 CAP_CHAIN.cap_chain1 CAP_CHAIN.cap_chain_inv1.O DC 0
V125 CAP_CHAIN.cap_chain_inv1.I CAP_CHAIN.I DC 0
V126 CAP_CHAIN.cap_chain2 CAP_CHAIN.cap_chain_inv2.O DC 0
V127 CAP_CHAIN.cap_chain_inv2.I CAP_CHAIN.cap_chain1 DC 0
V128 CAP_CHAIN.cap_chain3 CAP_CHAIN.cap_chain_inv3.O DC 0
V129 CAP_CHAIN.cap_chain_inv3.I CAP_CHAIN.cap_chain2 DC 0
V130 CAP_CHAIN.cap_chain4 CAP_CHAIN.cap_chain_inv4.O DC 0
V131 CAP_CHAIN.cap_chain_inv4.I CAP_CHAIN.cap_chain3 DC 0
V132 CAP_CHAIN.cap_chain5 CAP_CHAIN.cap_chain_inv5.O DC 0
V133 CAP_CHAIN.cap_chain_inv5.I CAP_CHAIN.cap_chain4 DC 0
V134 CAP_CHAIN.cap_chain6 CAP_CHAIN.cap_chain_inv6.O DC 0
V135 CAP_CHAIN.cap_chain_inv6.I CAP_CHAIN.cap_chain5 DC 0
V136 CAP_CHAIN.cap_chain7 CAP_CHAIN.cap_chain_inv7.O DC 0
V137 CAP_CHAIN.cap_chain_inv7.I CAP_CHAIN.cap_chain6 DC 0
V138 CAP_CHAIN.cap_chain8 CAP_CHAIN.cap_chain_inv8.O DC 0
V139 CAP_CHAIN.cap_chain_inv8.I CAP_CHAIN.cap_chain7 DC 0
V140 CAP_CHAIN.cap_chain9 CAP_CHAIN.cap_chain_inv9.O DC 0
V141 CAP_CHAIN.cap_chain_inv9.I CAP_CHAIN.cap_chain8 DC 0
V142 CAP_CHAIN.cap_chain10 CAP_CHAIN.cap_chain_inv10.O DC 0
V143 CAP_CHAIN.cap_chain_inv10.I CAP_CHAIN.cap_chain9 DC 0
V144 FINISH_CHAIN.finish_chain1 FINISH_CHAIN.finish_chain_inv1.O DC 0
V145 FINISH_CHAIN.finish_chain_inv1.I FINISH_CHAIN.I DC 0
V146 FINISH_CHAIN.finish_chain2 FINISH_CHAIN.finish_chain_inv2.O DC 0
V147 FINISH_CHAIN.finish_chain_inv2.I FINISH_CHAIN.finish_chain1 DC 0
V148 FINISH_CHAIN.finish_chain3 FINISH_CHAIN.finish_chain_inv3.O DC 0
V149 FINISH_CHAIN.finish_chain_inv3.I FINISH_CHAIN.finish_chain2 DC 0
V150 FINISH_CHAIN.finish_chain4 FINISH_CHAIN.finish_chain_inv4.O DC 0
V151 FINISH_CHAIN.finish_chain_inv4.I FINISH_CHAIN.finish_chain3 DC 0
V152 FINISH_CHAIN.finish_chain5 FINISH_CHAIN.finish_chain_inv5.O DC 0
V153 FINISH_CHAIN.finish_chain_inv5.I FINISH_CHAIN.finish_chain4 DC 0
V154 FINISH_CHAIN.finish_chain6 FINISH_CHAIN.finish_chain_inv6.O DC 0
V155 FINISH_CHAIN.finish_chain_inv6.I FINISH_CHAIN.finish_chain5 DC 0
V156 FINISH_CHAIN.finish_chain7 FINISH_CHAIN.finish_chain_inv7.O DC 0
V157 FINISH_CHAIN.finish_chain_inv7.I FINISH_CHAIN.finish_chain6 DC 0
V158 FINISH_CHAIN.finish_chain8 FINISH_CHAIN.finish_chain_inv8.O DC 0
V159 FINISH_CHAIN.finish_chain_inv8.I FINISH_CHAIN.finish_chain7 DC 0
V160 FINISH_CHAIN.finish_chain9 FINISH_CHAIN.finish_chain_inv9.O DC 0
V161 FINISH_CHAIN.finish_chain_inv9.I FINISH_CHAIN.finish_chain8 DC 0
V162 FINISH_CHAIN.finish_chain10 FINISH_CHAIN.finish_chain_inv10.O DC 0
V163 FINISH_CHAIN.finish_chain_inv10.I FINISH_CHAIN.finish_chain9 DC 0
V164 FINISH_CHAIN.finish_chain11 FINISH_CHAIN.finish_chain_inv11.O DC 0
V165 FINISH_CHAIN.finish_chain_inv11.I FINISH_CHAIN.finish_chain10 DC 0
V166 FINISH_CHAIN.finish_chain12 FINISH_CHAIN.finish_chain_inv12.O DC 0
V167 FINISH_CHAIN.finish_chain_inv12.I FINISH_CHAIN.finish_chain11 DC 0
V168 FINISH_CHAIN.finish_chain13 FINISH_CHAIN.finish_chain_inv13.O DC 0
V169 FINISH_CHAIN.finish_chain_inv13.I FINISH_CHAIN.finish_chain12 DC 0
V170 FINISH_CHAIN.finish_chain14 FINISH_CHAIN.finish_chain_inv14.O DC 0
V171 FINISH_CHAIN.finish_chain_inv14.I FINISH_CHAIN.finish_chain13 DC 0
V172 FINISH_CHAIN.Ob FINISH_CHAIN.finish_chain_inv15.O DC 0
V173 FINISH_CHAIN.finish_chain_inv15.I FINISH_CHAIN.finish_chain14 DC 0
V174 FINISH_CHAIN.O FINISH_CHAIN.finish_chain_inv16.O DC 0
V175 FINISH_CHAIN.finish_chain_inv16.I FINISH_CHAIN.Ob DC 0
V176 FALLING_COMP.Db_Minus FALLING_COMP.INV_DM.O DC 0
V177 FALLING_COMP.INV_DM.I FALLING_COMP.D_Minus DC 0
V178 CAP_CHAIN.cap_chain11 CAP_CHAIN.cap_chain_inv11.O DC 0
V179 CAP_CHAIN.cap_chain_inv11.I CAP_CHAIN.cap_chain10 DC 0
V180 CAP_CHAIN.cap_chain12 CAP_CHAIN.cap_chain_inv12.O DC 0
V181 CAP_CHAIN.cap_chain_inv12.I CAP_CHAIN.cap_chain11 DC 0
V182 CAP_CHAIN.cap_chain13 CAP_CHAIN.cap_chain_inv13.O DC 0
V183 CAP_CHAIN.cap_chain_inv13.I CAP_CHAIN.cap_chain12 DC 0
V184 CAP_CHAIN.cap_chain14 CAP_CHAIN.cap_chain_inv14.O DC 0
V185 CAP_CHAIN.cap_chain_inv14.I CAP_CHAIN.cap_chain13 DC 0
V186 CAP_CHAIN.cap_chain15 CAP_CHAIN.cap_chain_inv15.O DC 0
V187 CAP_CHAIN.cap_chain_inv15.I CAP_CHAIN.cap_chain14 DC 0
V188 CAP_CHAIN.O CAP_CHAIN.cap_chain_inv16.O DC 0
V189 CAP_CHAIN.cap_chain_inv16.I CAP_CHAIN.cap_chain15 DC 0
V190 FALLING_COMP.Db_Plus FALLING_COMP.INV_DP.O DC 0
V191 FALLING_COMP.INV_DP.I FALLING_COMP.D_Plus DC 0
V192 FALLING_COMP.Qb FALLING_COMP.SR_MEM.Qb DC 0
V193 FALLING_COMP.Q FALLING_COMP.SR_MEM.Q DC 0
V194 FALLING_COMP.SR_MEM.Rb FALLING_COMP.Db_Minus DC 0
V195 FALLING_COMP.SR_MEM.Sb FALLING_COMP.Db_Plus DC 0
V196 FALLING_COMP.Qb_b FALLING_COMP.INV_Qb.O DC 0
V197 FALLING_COMP.INV_Qb.I FALLING_COMP.Qb DC 0
V198 FALLING_COMP.Done FALLING_COMP.NAND2_COMP.O DC 0
V199 FALLING_COMP.NAND2_COMP.B FALLING_COMP.D_Minus DC 0
V200 FALLING_COMP.NAND2_COMP.A FALLING_COMP.D_Plus DC 0
V201 CLOCK_GEN.FinishB_Delay CLOCK_GEN.INV_F.O DC 0
V202 CLOCK_GEN.INV_F.I CLOCK_GEN.Finish_Delay DC 0
V203 CLOCK_GEN.Set_OE CLOCK_GEN.NAND_DF.O DC 0
V204 CLOCK_GEN.NAND_DF.B CLOCK_GEN.FinishB_Delay DC 0
V205 CLOCK_GEN.NAND_DF.A CLOCK_GEN.Done_Falling DC 0
V206 RISING_COMP.Done RISING_COMP.NAND2_COMP.O DC 0
V207 RISING_COMP.NAND2_COMP.B RISING_COMP.D_Minus DC 0
V208 RISING_COMP.NAND2_COMP.A RISING_COMP.D_Plus DC 0
V209 CLOCK_GEN.Reset_OE CLOCK_GEN.NAND_DR.O DC 0
V210 CLOCK_GEN.NAND_DR.B CLOCK_GEN.Finish_Delay DC 0
V211 CLOCK_GEN.NAND_DR.A CLOCK_GEN.Done_Rising DC 0
V212 CLOCK_GEN.OE_Falling CLOCK_GEN.SR_OE.Q DC 0
V213 CLOCK_GEN.SR_OE.Rb CLOCK_GEN.Reset_OE DC 0
V214 CLOCK_GEN.SR_OE.Sb CLOCK_GEN.Set_OE DC 0
V215 FALLING_COMP.Y FALLING_COMP.NAND3_COMP.O DC 0
V216 FALLING_COMP.NAND3_COMP.C FALLING_COMP.Output_Enable DC 0
V217 FALLING_COMP.NAND3_COMP.B FALLING_COMP.Db_Plus DC 0
V218 FALLING_COMP.NAND3_COMP.A FALLING_COMP.Qb_b DC 0
V219 FALLING_COUNTER.D.0 FALLING_COUNTER.COUNT_SUB_INV0.O DC 0
V220 FALLING_COUNTER.COUNT_SUB_INV0.I FALLING_COUNTER.O.0 DC 0
V221 FALLING_COUNTER.O.0 FALLING_COUNTER.COUNT_SUB_DFF0.Q DC 0
V222 FALLING_COUNTER.COUNT_SUB_DFF0.RSTb FALLING_COUNTER.RSTb DC 0
V223 FALLING_COUNTER.COUNT_SUB_DFF0.D FALLING_COUNTER.D.0 DC 0
V224 FALLING_COUNTER.COUNT_SUB_DFF0.CLK FALLING_COUNTER.CLK DC 0
V225 FALLING_COUNTER.D.1 FALLING_COUNTER.COUNT_SUB_INV1.O DC 0
V226 FALLING_COUNTER.COUNT_SUB_INV1.I FALLING_COUNTER.O.1 DC 0
V227 FALLING_COUNTER.O.1 FALLING_COUNTER.COUNT_SUB_DFF1.Q DC 0
V228 FALLING_COUNTER.COUNT_SUB_DFF1.RSTb FALLING_COUNTER.RSTb DC 0
V229 FALLING_COUNTER.COUNT_SUB_DFF1.D FALLING_COUNTER.D.1 DC 0
V230 FALLING_COUNTER.COUNT_SUB_DFF1.CLK FALLING_COUNTER.O.0 DC 0
V231 FALLING_COUNTER.D.2 FALLING_COUNTER.COUNT_SUB_INV2.O DC 0
V232 FALLING_COUNTER.COUNT_SUB_INV2.I FALLING_COUNTER.O.2 DC 0
V233 FALLING_COUNTER.O.2 FALLING_COUNTER.COUNT_SUB_DFF2.Q DC 0
V234 FALLING_COUNTER.COUNT_SUB_DFF2.RSTb FALLING_COUNTER.RSTb DC 0
V235 FALLING_COUNTER.COUNT_SUB_DFF2.D FALLING_COUNTER.D.2 DC 0
V236 FALLING_COUNTER.COUNT_SUB_DFF2.CLK FALLING_COUNTER.O.1 DC 0
V237 FALLING_COUNTER.D.3 FALLING_COUNTER.COUNT_SUB_INV3.O DC 0
V238 FALLING_COUNTER.COUNT_SUB_INV3.I FALLING_COUNTER.O.3 DC 0
V239 FALLING_COUNTER.O.3 FALLING_COUNTER.COUNT_SUB_DFF3.Q DC 0
V240 FALLING_COUNTER.COUNT_SUB_DFF3.RSTb FALLING_COUNTER.RSTb DC 0
V241 FALLING_COUNTER.COUNT_SUB_DFF3.D FALLING_COUNTER.D.3 DC 0
V242 FALLING_COUNTER.COUNT_SUB_DFF3.CLK FALLING_COUNTER.O.2 DC 0
V243 FALLING_COUNTER.D.4 FALLING_COUNTER.COUNT_SUB_INV4.O DC 0
V244 FALLING_COUNTER.COUNT_SUB_INV4.I FALLING_COUNTER.O.4 DC 0
V245 FALLING_COUNTER.O.4 FALLING_COUNTER.COUNT_SUB_DFF4.Q DC 0
V246 FALLING_COUNTER.COUNT_SUB_DFF4.RSTb FALLING_COUNTER.RSTb DC 0
V247 FALLING_COUNTER.COUNT_SUB_DFF4.D FALLING_COUNTER.D.4 DC 0
V248 FALLING_COUNTER.COUNT_SUB_DFF4.CLK FALLING_COUNTER.O.3 DC 0
V249 FALLING_COUNTER.D.5 FALLING_COUNTER.COUNT_SUB_INV5.O DC 0
V250 FALLING_COUNTER.COUNT_SUB_INV5.I FALLING_COUNTER.O.5 DC 0
V251 FALLING_COUNTER.O.5 FALLING_COUNTER.COUNT_SUB_DFF5.Q DC 0
V252 FALLING_COUNTER.COUNT_SUB_DFF5.RSTb FALLING_COUNTER.RSTb DC 0
V253 FALLING_COUNTER.COUNT_SUB_DFF5.D FALLING_COUNTER.D.5 DC 0
V254 FALLING_COUNTER.COUNT_SUB_DFF5.CLK FALLING_COUNTER.O.4 DC 0
V255 FALLING_COUNTER.D.6 FALLING_COUNTER.COUNT_SUB_INV6.O DC 0
V256 FALLING_COUNTER.COUNT_SUB_INV6.I FALLING_COUNTER.O.6 DC 0
V257 FALLING_COUNTER.O.6 FALLING_COUNTER.COUNT_SUB_DFF6.Q DC 0
V258 FALLING_COUNTER.COUNT_SUB_DFF6.RSTb FALLING_COUNTER.RSTb DC 0
V259 FALLING_COUNTER.COUNT_SUB_DFF6.D FALLING_COUNTER.D.6 DC 0
V260 FALLING_COUNTER.COUNT_SUB_DFF6.CLK FALLING_COUNTER.O.5 DC 0
V261 FALLING_COUNTER.D.7 FALLING_COUNTER.COUNT_SUB_INV7.O DC 0
V262 FALLING_COUNTER.COUNT_SUB_INV7.I FALLING_COUNTER.O.7 DC 0
V263 FALLING_COUNTER.O.7 FALLING_COUNTER.COUNT_SUB_DFF7.Q DC 0
V264 FALLING_COUNTER.COUNT_SUB_DFF7.RSTb FALLING_COUNTER.RSTb DC 0
V265 FALLING_COUNTER.COUNT_SUB_DFF7.D FALLING_COUNTER.D.7 DC 0
V266 FALLING_COUNTER.COUNT_SUB_DFF7.CLK FALLING_COUNTER.O.6 DC 0
V267 FALLING_COUNTER.D.8 FALLING_COUNTER.COUNT_SUB_INV8.O DC 0
V268 FALLING_COUNTER.COUNT_SUB_INV8.I FALLING_COUNTER.O.8 DC 0
V269 FALLING_COUNTER.O.8 FALLING_COUNTER.COUNT_SUB_DFF8.Q DC 0
V270 FALLING_COUNTER.COUNT_SUB_DFF8.RSTb FALLING_COUNTER.RSTb DC 0
V271 FALLING_COUNTER.COUNT_SUB_DFF8.D FALLING_COUNTER.D.8 DC 0
V272 FALLING_COUNTER.COUNT_SUB_DFF8.CLK FALLING_COUNTER.O.7 DC 0
V273 FALLING_COUNTER.D.9 FALLING_COUNTER.COUNT_SUB_INV9.O DC 0
V274 FALLING_COUNTER.COUNT_SUB_INV9.I FALLING_COUNTER.O.9 DC 0
V275 FALLING_COUNTER.O.9 FALLING_COUNTER.COUNT_SUB_DFF9.Q DC 0
V276 FALLING_COUNTER.COUNT_SUB_DFF9.RSTb FALLING_COUNTER.RSTb DC 0
V277 FALLING_COUNTER.COUNT_SUB_DFF9.D FALLING_COUNTER.D.9 DC 0
V278 FALLING_COUNTER.COUNT_SUB_DFF9.CLK FALLING_COUNTER.O.8 DC 0
V279 FALLING_COUNTER.D.10 FALLING_COUNTER.COUNT_SUB_INV10.O DC 0
V280 FALLING_COUNTER.COUNT_SUB_INV10.I FALLING_COUNTER.O.10 DC 0
V281 FALLING_COUNTER.O.10 FALLING_COUNTER.COUNT_SUB_DFF10.Q DC 0
V282 FALLING_COUNTER.COUNT_SUB_DFF10.RSTb FALLING_COUNTER.RSTb DC 0
V283 FALLING_COUNTER.COUNT_SUB_DFF10.D FALLING_COUNTER.D.10 DC 0
V284 FALLING_COUNTER.COUNT_SUB_DFF10.CLK FALLING_COUNTER.O.9 DC 0
V285 FALLING_COUNTER.D.11 FALLING_COUNTER.COUNT_SUB_INV11.O DC 0
V286 FALLING_COUNTER.COUNT_SUB_INV11.I FALLING_COUNTER.O.11 DC 0
V287 FALLING_COUNTER.O.11 FALLING_COUNTER.COUNT_SUB_DFF11.Q DC 0
V288 FALLING_COUNTER.COUNT_SUB_DFF11.RSTb FALLING_COUNTER.RSTb DC 0
V289 FALLING_COUNTER.COUNT_SUB_DFF11.D FALLING_COUNTER.D.11 DC 0
V290 FALLING_COUNTER.COUNT_SUB_DFF11.CLK FALLING_COUNTER.O.10 DC 0
V291 FALLING_COUNTER.D.12 FALLING_COUNTER.COUNT_SUB_INV12.O DC 0
V292 FALLING_COUNTER.COUNT_SUB_INV12.I FALLING_COUNTER.O.12 DC 0
V293 FALLING_COUNTER.O.12 FALLING_COUNTER.COUNT_SUB_DFF12.Q DC 0
V294 FALLING_COUNTER.COUNT_SUB_DFF12.RSTb FALLING_COUNTER.RSTb DC 0
V295 FALLING_COUNTER.COUNT_SUB_DFF12.D FALLING_COUNTER.D.12 DC 0
V296 FALLING_COUNTER.COUNT_SUB_DFF12.CLK FALLING_COUNTER.O.11 DC 0
V297 FALLING_COUNTER.D.13 FALLING_COUNTER.COUNT_SUB_INV13.O DC 0
V298 FALLING_COUNTER.COUNT_SUB_INV13.I FALLING_COUNTER.O.13 DC 0
V299 FALLING_COUNTER.O.13 FALLING_COUNTER.COUNT_SUB_DFF13.Q DC 0
V300 FALLING_COUNTER.COUNT_SUB_DFF13.RSTb FALLING_COUNTER.RSTb DC 0
V301 FALLING_COUNTER.COUNT_SUB_DFF13.D FALLING_COUNTER.D.13 DC 0
V302 FALLING_COUNTER.COUNT_SUB_DFF13.CLK FALLING_COUNTER.O.12 DC 0
V303 FALLING_COUNTER.D.14 FALLING_COUNTER.COUNT_SUB_INV14.O DC 0
V304 FALLING_COUNTER.COUNT_SUB_INV14.I FALLING_COUNTER.O.14 DC 0
V305 FALLING_COUNTER.O.14 FALLING_COUNTER.COUNT_SUB_DFF14.Q DC 0
V306 FALLING_COUNTER.COUNT_SUB_DFF14.RSTb FALLING_COUNTER.RSTb DC 0
V307 FALLING_COUNTER.COUNT_SUB_DFF14.D FALLING_COUNTER.D.14 DC 0
V308 FALLING_COUNTER.COUNT_SUB_DFF14.CLK FALLING_COUNTER.O.13 DC 0
V309 FALLING_COMP.Q_b FALLING_COMP.INV_Q.O DC 0
V310 FALLING_COMP.INV_Q.I FALLING_COMP.Q DC 0
V311 RISING_COMP.Db_Plus RISING_COMP.INV_DP.O DC 0
V312 RISING_COMP.INV_DP.I RISING_COMP.D_Plus DC 0
V313 RISING_COMP.Db_Minus RISING_COMP.INV_DM.O DC 0
V314 RISING_COMP.INV_DM.I RISING_COMP.D_Minus DC 0
V315 RISING_COMP.Qb RISING_COMP.SR_MEM.Qb DC 0
V316 RISING_COMP.Q RISING_COMP.SR_MEM.Q DC 0
V317 RISING_COMP.SR_MEM.Rb RISING_COMP.Db_Minus DC 0
V318 RISING_COMP.SR_MEM.Sb RISING_COMP.Db_Plus DC 0
V319 RISING_COMP.Qb_b RISING_COMP.INV_Qb.O DC 0
V320 RISING_COMP.INV_Qb.I RISING_COMP.Qb DC 0
V321 CLOCK_GEN.OE_Rising CLOCK_GEN.INV_OE.O DC 0
V322 CLOCK_GEN.INV_OE.I CLOCK_GEN.OE_Falling DC 0
V323 RISING_COMP.Y RISING_COMP.NAND3_COMP.O DC 0
V324 RISING_COMP.NAND3_COMP.C RISING_COMP.Output_Enable DC 0
V325 RISING_COMP.NAND3_COMP.B RISING_COMP.Db_Plus DC 0
V326 RISING_COMP.NAND3_COMP.A RISING_COMP.Qb_b DC 0
V327 RISING_COMP.Q_b RISING_COMP.INV_Q.O DC 0
V328 RISING_COMP.INV_Q.I RISING_COMP.Q DC 0
V329 FINISH_COMP.Db_Minus FINISH_COMP.INV_DM.O DC 0
V330 FINISH_COMP.INV_DM.I FINISH_COMP.D_Minus DC 0
V331 FINISH_COMP.Db_Plus FINISH_COMP.INV_DP.O DC 0
V332 FINISH_COMP.INV_DP.I FINISH_COMP.D_Plus DC 0
V333 FINISH_COMP.Qb FINISH_COMP.SR_MEM.Qb DC 0
V334 FINISH_COMP.Q FINISH_COMP.SR_MEM.Q DC 0
V335 FINISH_COMP.SR_MEM.Rb FINISH_COMP.Db_Minus DC 0
V336 FINISH_COMP.SR_MEM.Sb FINISH_COMP.Db_Plus DC 0
V337 FINISH_COMP.Qb_b FINISH_COMP.INV_Qb.O DC 0
V338 FINISH_COMP.INV_Qb.I FINISH_COMP.Qb DC 0
V339 FINISH_COMP.Y FINISH_COMP.NAND3_COMP.O DC 0
V340 FINISH_COMP.NAND3_COMP.C FINISH_COMP.Output_Enable DC 0
V341 FINISH_COMP.NAND3_COMP.B FINISH_COMP.Db_Plus DC 0
V342 FINISH_COMP.NAND3_COMP.A FINISH_COMP.Qb_b DC 0
V343 FINISH_COMP.Done FINISH_COMP.NAND2_COMP.O DC 0
V344 FINISH_COMP.NAND2_COMP.B FINISH_COMP.D_Minus DC 0
V345 FINISH_COMP.NAND2_COMP.A FINISH_COMP.D_Plus DC 0
V346 FINISH_COMP.Q_b FINISH_COMP.INV_Q.O DC 0
V347 FINISH_COMP.INV_Q.I FINISH_COMP.Q DC 0
V348 CLOCK_GEN.ResetB CLOCK_GEN.INV_R.O DC 0
V349 CLOCK_GEN.INV_R.I CLOCK_GEN.Reset DC 0
V350 CLOCK_GEN.Conv_Finish CLOCK_GEN.SR_Op.Q DC 0
V351 CLOCK_GEN.SR_Op.Rb CLOCK_GEN.ResetB DC 0
V352 CLOCK_GEN.SR_Op.Sb CLOCK_GEN.Finish DC 0
V353 CLOCK_GEN.Sense CLOCK_GEN.NOR_CLK.O DC 0
V354 CLOCK_GEN.NOR_CLK.B CLOCK_GEN.Conv_Finish DC 0
V355 CLOCK_GEN.NOR_CLK.A CLOCK_GEN.Reset DC 0
V356 CLOCK_GEN.CLKb CLOCK_GEN.NAND_CLK.O DC 0
V357 CLOCK_GEN.NAND_CLK.B CLOCK_GEN.Sense DC 0
V358 CLOCK_GEN.NAND_CLK.A CLOCK_GEN.OE_Falling DC 0
V359 CLOCK_GEN.Next_Edge CLOCK_GEN.NOT_CLK.O DC 0
V360 CLOCK_GEN.NOT_CLK.I CLOCK_GEN.CLKb DC 0
V361 RISING_COUNTER.D.0 RISING_COUNTER.COUNT_SUB_INV0.O DC 0
V362 RISING_COUNTER.COUNT_SUB_INV0.I RISING_COUNTER.O.0 DC 0
V363 RISING_COUNTER.O.0 RISING_COUNTER.COUNT_SUB_DFF0.Q DC 0
V364 RISING_COUNTER.COUNT_SUB_DFF0.RSTb RISING_COUNTER.RSTb DC 0
V365 RISING_COUNTER.COUNT_SUB_DFF0.D RISING_COUNTER.D.0 DC 0
V366 RISING_COUNTER.COUNT_SUB_DFF0.CLK RISING_COUNTER.CLK DC 0
V367 RISING_COUNTER.D.1 RISING_COUNTER.COUNT_SUB_INV1.O DC 0
V368 RISING_COUNTER.COUNT_SUB_INV1.I RISING_COUNTER.O.1 DC 0
V369 RISING_COUNTER.O.1 RISING_COUNTER.COUNT_SUB_DFF1.Q DC 0
V370 RISING_COUNTER.COUNT_SUB_DFF1.RSTb RISING_COUNTER.RSTb DC 0
V371 RISING_COUNTER.COUNT_SUB_DFF1.D RISING_COUNTER.D.1 DC 0
V372 RISING_COUNTER.COUNT_SUB_DFF1.CLK RISING_COUNTER.O.0 DC 0
V373 RISING_COUNTER.D.2 RISING_COUNTER.COUNT_SUB_INV2.O DC 0
V374 RISING_COUNTER.COUNT_SUB_INV2.I RISING_COUNTER.O.2 DC 0
V375 RISING_COUNTER.O.2 RISING_COUNTER.COUNT_SUB_DFF2.Q DC 0
V376 RISING_COUNTER.COUNT_SUB_DFF2.RSTb RISING_COUNTER.RSTb DC 0
V377 RISING_COUNTER.COUNT_SUB_DFF2.D RISING_COUNTER.D.2 DC 0
V378 RISING_COUNTER.COUNT_SUB_DFF2.CLK RISING_COUNTER.O.1 DC 0
V379 RISING_COUNTER.D.3 RISING_COUNTER.COUNT_SUB_INV3.O DC 0
V380 RISING_COUNTER.COUNT_SUB_INV3.I RISING_COUNTER.O.3 DC 0
V381 RISING_COUNTER.O.3 RISING_COUNTER.COUNT_SUB_DFF3.Q DC 0
V382 RISING_COUNTER.COUNT_SUB_DFF3.RSTb RISING_COUNTER.RSTb DC 0
V383 RISING_COUNTER.COUNT_SUB_DFF3.D RISING_COUNTER.D.3 DC 0
V384 RISING_COUNTER.COUNT_SUB_DFF3.CLK RISING_COUNTER.O.2 DC 0
V385 RISING_COUNTER.D.4 RISING_COUNTER.COUNT_SUB_INV4.O DC 0
V386 RISING_COUNTER.COUNT_SUB_INV4.I RISING_COUNTER.O.4 DC 0
V387 RISING_COUNTER.O.4 RISING_COUNTER.COUNT_SUB_DFF4.Q DC 0
V388 RISING_COUNTER.COUNT_SUB_DFF4.RSTb RISING_COUNTER.RSTb DC 0
V389 RISING_COUNTER.COUNT_SUB_DFF4.D RISING_COUNTER.D.4 DC 0
V390 RISING_COUNTER.COUNT_SUB_DFF4.CLK RISING_COUNTER.O.3 DC 0
V391 RISING_COUNTER.D.5 RISING_COUNTER.COUNT_SUB_INV5.O DC 0
V392 RISING_COUNTER.COUNT_SUB_INV5.I RISING_COUNTER.O.5 DC 0
V393 RISING_COUNTER.O.5 RISING_COUNTER.COUNT_SUB_DFF5.Q DC 0
V394 RISING_COUNTER.COUNT_SUB_DFF5.RSTb RISING_COUNTER.RSTb DC 0
V395 RISING_COUNTER.COUNT_SUB_DFF5.D RISING_COUNTER.D.5 DC 0
V396 RISING_COUNTER.COUNT_SUB_DFF5.CLK RISING_COUNTER.O.4 DC 0
V397 RISING_COUNTER.D.6 RISING_COUNTER.COUNT_SUB_INV6.O DC 0
V398 RISING_COUNTER.COUNT_SUB_INV6.I RISING_COUNTER.O.6 DC 0
V399 RISING_COUNTER.O.6 RISING_COUNTER.COUNT_SUB_DFF6.Q DC 0
V400 RISING_COUNTER.COUNT_SUB_DFF6.RSTb RISING_COUNTER.RSTb DC 0
V401 RISING_COUNTER.COUNT_SUB_DFF6.D RISING_COUNTER.D.6 DC 0
V402 RISING_COUNTER.COUNT_SUB_DFF6.CLK RISING_COUNTER.O.5 DC 0
V403 RISING_COUNTER.D.7 RISING_COUNTER.COUNT_SUB_INV7.O DC 0
V404 RISING_COUNTER.COUNT_SUB_INV7.I RISING_COUNTER.O.7 DC 0
V405 RISING_COUNTER.O.7 RISING_COUNTER.COUNT_SUB_DFF7.Q DC 0
V406 RISING_COUNTER.COUNT_SUB_DFF7.RSTb RISING_COUNTER.RSTb DC 0
V407 RISING_COUNTER.COUNT_SUB_DFF7.D RISING_COUNTER.D.7 DC 0
V408 RISING_COUNTER.COUNT_SUB_DFF7.CLK RISING_COUNTER.O.6 DC 0
V409 RISING_COUNTER.D.8 RISING_COUNTER.COUNT_SUB_INV8.O DC 0
V410 RISING_COUNTER.COUNT_SUB_INV8.I RISING_COUNTER.O.8 DC 0
V411 RISING_COUNTER.O.8 RISING_COUNTER.COUNT_SUB_DFF8.Q DC 0
V412 RISING_COUNTER.COUNT_SUB_DFF8.RSTb RISING_COUNTER.RSTb DC 0
V413 RISING_COUNTER.COUNT_SUB_DFF8.D RISING_COUNTER.D.8 DC 0
V414 RISING_COUNTER.COUNT_SUB_DFF8.CLK RISING_COUNTER.O.7 DC 0
V415 RISING_COUNTER.D.9 RISING_COUNTER.COUNT_SUB_INV9.O DC 0
V416 RISING_COUNTER.COUNT_SUB_INV9.I RISING_COUNTER.O.9 DC 0
V417 RISING_COUNTER.O.9 RISING_COUNTER.COUNT_SUB_DFF9.Q DC 0
V418 RISING_COUNTER.COUNT_SUB_DFF9.RSTb RISING_COUNTER.RSTb DC 0
V419 RISING_COUNTER.COUNT_SUB_DFF9.D RISING_COUNTER.D.9 DC 0
V420 RISING_COUNTER.COUNT_SUB_DFF9.CLK RISING_COUNTER.O.8 DC 0
V421 RISING_COUNTER.D.10 RISING_COUNTER.COUNT_SUB_INV10.O DC 0
V422 RISING_COUNTER.COUNT_SUB_INV10.I RISING_COUNTER.O.10 DC 0
V423 RISING_COUNTER.O.10 RISING_COUNTER.COUNT_SUB_DFF10.Q DC 0
V424 RISING_COUNTER.COUNT_SUB_DFF10.RSTb RISING_COUNTER.RSTb DC 0
V425 RISING_COUNTER.COUNT_SUB_DFF10.D RISING_COUNTER.D.10 DC 0
V426 RISING_COUNTER.COUNT_SUB_DFF10.CLK RISING_COUNTER.O.9 DC 0
V427 RISING_COUNTER.D.11 RISING_COUNTER.COUNT_SUB_INV11.O DC 0
V428 RISING_COUNTER.COUNT_SUB_INV11.I RISING_COUNTER.O.11 DC 0
V429 RISING_COUNTER.O.11 RISING_COUNTER.COUNT_SUB_DFF11.Q DC 0
V430 RISING_COUNTER.COUNT_SUB_DFF11.RSTb RISING_COUNTER.RSTb DC 0
V431 RISING_COUNTER.COUNT_SUB_DFF11.D RISING_COUNTER.D.11 DC 0
V432 RISING_COUNTER.COUNT_SUB_DFF11.CLK RISING_COUNTER.O.10 DC 0
V433 RISING_COUNTER.D.12 RISING_COUNTER.COUNT_SUB_INV12.O DC 0
V434 RISING_COUNTER.COUNT_SUB_INV12.I RISING_COUNTER.O.12 DC 0
V435 RISING_COUNTER.O.12 RISING_COUNTER.COUNT_SUB_DFF12.Q DC 0
V436 RISING_COUNTER.COUNT_SUB_DFF12.RSTb RISING_COUNTER.RSTb DC 0
V437 RISING_COUNTER.COUNT_SUB_DFF12.D RISING_COUNTER.D.12 DC 0
V438 RISING_COUNTER.COUNT_SUB_DFF12.CLK RISING_COUNTER.O.11 DC 0
V439 RISING_COUNTER.D.13 RISING_COUNTER.COUNT_SUB_INV13.O DC 0
V440 RISING_COUNTER.COUNT_SUB_INV13.I RISING_COUNTER.O.13 DC 0
V441 RISING_COUNTER.O.13 RISING_COUNTER.COUNT_SUB_DFF13.Q DC 0
V442 RISING_COUNTER.COUNT_SUB_DFF13.RSTb RISING_COUNTER.RSTb DC 0
V443 RISING_COUNTER.COUNT_SUB_DFF13.D RISING_COUNTER.D.13 DC 0
V444 RISING_COUNTER.COUNT_SUB_DFF13.CLK RISING_COUNTER.O.12 DC 0
V445 RISING_COUNTER.D.14 RISING_COUNTER.COUNT_SUB_INV14.O DC 0
V446 RISING_COUNTER.COUNT_SUB_INV14.I RISING_COUNTER.O.14 DC 0
V447 RISING_COUNTER.O.14 RISING_COUNTER.COUNT_SUB_DFF14.Q DC 0
V448 RISING_COUNTER.COUNT_SUB_DFF14.RSTb RISING_COUNTER.RSTb DC 0
V449 RISING_COUNTER.COUNT_SUB_DFF14.D RISING_COUNTER.D.14 DC 0
V450 RISING_COUNTER.COUNT_SUB_DFF14.CLK RISING_COUNTER.O.13 DC 0
V451 FALLING_COUNTER.D.15 FALLING_COUNTER.COUNT_SUB_INV15.O DC 0
V452 FALLING_COUNTER.COUNT_SUB_INV15.I FALLING_COUNTER.O.15 DC 0
V453 FALLING_COUNTER.O.15 FALLING_COUNTER.COUNT_SUB_DFF15.Q DC 0
V454 FALLING_COUNTER.COUNT_SUB_DFF15.RSTb FALLING_COUNTER.RSTb DC 0
V455 FALLING_COUNTER.COUNT_SUB_DFF15.D FALLING_COUNTER.D.15 DC 0
V456 FALLING_COUNTER.COUNT_SUB_DFF15.CLK FALLING_COUNTER.O.14 DC 0
V457 FULL_COUNTER.D.0 FULL_COUNTER.COUNT_SUB_INV0.O DC 0
V458 FULL_COUNTER.COUNT_SUB_INV0.I FULL_COUNTER.O.0 DC 0
V459 FULL_COUNTER.O.0 FULL_COUNTER.COUNT_SUB_DFF0.Q DC 0
V460 FULL_COUNTER.COUNT_SUB_DFF0.RSTb FULL_COUNTER.RSTb DC 0
V461 FULL_COUNTER.COUNT_SUB_DFF0.D FULL_COUNTER.D.0 DC 0
V462 FULL_COUNTER.COUNT_SUB_DFF0.CLK FULL_COUNTER.CLK DC 0
V463 FULL_COUNTER.D.1 FULL_COUNTER.COUNT_SUB_INV1.O DC 0
V464 FULL_COUNTER.COUNT_SUB_INV1.I FULL_COUNTER.O.1 DC 0
V465 FULL_COUNTER.O.1 FULL_COUNTER.COUNT_SUB_DFF1.Q DC 0
V466 FULL_COUNTER.COUNT_SUB_DFF1.RSTb FULL_COUNTER.RSTb DC 0
V467 FULL_COUNTER.COUNT_SUB_DFF1.D FULL_COUNTER.D.1 DC 0
V468 FULL_COUNTER.COUNT_SUB_DFF1.CLK FULL_COUNTER.O.0 DC 0
V469 FULL_COUNTER.D.2 FULL_COUNTER.COUNT_SUB_INV2.O DC 0
V470 FULL_COUNTER.COUNT_SUB_INV2.I FULL_COUNTER.O.2 DC 0
V471 FULL_COUNTER.O.2 FULL_COUNTER.COUNT_SUB_DFF2.Q DC 0
V472 FULL_COUNTER.COUNT_SUB_DFF2.RSTb FULL_COUNTER.RSTb DC 0
V473 FULL_COUNTER.COUNT_SUB_DFF2.D FULL_COUNTER.D.2 DC 0
V474 FULL_COUNTER.COUNT_SUB_DFF2.CLK FULL_COUNTER.O.1 DC 0
V475 FULL_COUNTER.D.3 FULL_COUNTER.COUNT_SUB_INV3.O DC 0
V476 FULL_COUNTER.COUNT_SUB_INV3.I FULL_COUNTER.O.3 DC 0
V477 FULL_COUNTER.O.3 FULL_COUNTER.COUNT_SUB_DFF3.Q DC 0
V478 FULL_COUNTER.COUNT_SUB_DFF3.RSTb FULL_COUNTER.RSTb DC 0
V479 FULL_COUNTER.COUNT_SUB_DFF3.D FULL_COUNTER.D.3 DC 0
V480 FULL_COUNTER.COUNT_SUB_DFF3.CLK FULL_COUNTER.O.2 DC 0
V481 FULL_COUNTER.D.4 FULL_COUNTER.COUNT_SUB_INV4.O DC 0
V482 FULL_COUNTER.COUNT_SUB_INV4.I FULL_COUNTER.O.4 DC 0
V483 FULL_COUNTER.O.4 FULL_COUNTER.COUNT_SUB_DFF4.Q DC 0
V484 FULL_COUNTER.COUNT_SUB_DFF4.RSTb FULL_COUNTER.RSTb DC 0
V485 FULL_COUNTER.COUNT_SUB_DFF4.D FULL_COUNTER.D.4 DC 0
V486 FULL_COUNTER.COUNT_SUB_DFF4.CLK FULL_COUNTER.O.3 DC 0
V487 FULL_COUNTER.D.5 FULL_COUNTER.COUNT_SUB_INV5.O DC 0
V488 FULL_COUNTER.COUNT_SUB_INV5.I FULL_COUNTER.O.5 DC 0
V489 FULL_COUNTER.O.5 FULL_COUNTER.COUNT_SUB_DFF5.Q DC 0
V490 FULL_COUNTER.COUNT_SUB_DFF5.RSTb FULL_COUNTER.RSTb DC 0
V491 FULL_COUNTER.COUNT_SUB_DFF5.D FULL_COUNTER.D.5 DC 0
V492 FULL_COUNTER.COUNT_SUB_DFF5.CLK FULL_COUNTER.O.4 DC 0
V493 FULL_COUNTER.D.6 FULL_COUNTER.COUNT_SUB_INV6.O DC 0
V494 FULL_COUNTER.COUNT_SUB_INV6.I FULL_COUNTER.O.6 DC 0
V495 FULL_COUNTER.O.6 FULL_COUNTER.COUNT_SUB_DFF6.Q DC 0
V496 FULL_COUNTER.COUNT_SUB_DFF6.RSTb FULL_COUNTER.RSTb DC 0
V497 FULL_COUNTER.COUNT_SUB_DFF6.D FULL_COUNTER.D.6 DC 0
V498 FULL_COUNTER.COUNT_SUB_DFF6.CLK FULL_COUNTER.O.5 DC 0
V499 FULL_COUNTER.D.7 FULL_COUNTER.COUNT_SUB_INV7.O DC 0
V500 FULL_COUNTER.COUNT_SUB_INV7.I FULL_COUNTER.O.7 DC 0
V501 FULL_COUNTER.O.7 FULL_COUNTER.COUNT_SUB_DFF7.Q DC 0
V502 FULL_COUNTER.COUNT_SUB_DFF7.RSTb FULL_COUNTER.RSTb DC 0
V503 FULL_COUNTER.COUNT_SUB_DFF7.D FULL_COUNTER.D.7 DC 0
V504 FULL_COUNTER.COUNT_SUB_DFF7.CLK FULL_COUNTER.O.6 DC 0
V505 FULL_COUNTER.D.8 FULL_COUNTER.COUNT_SUB_INV8.O DC 0
V506 FULL_COUNTER.COUNT_SUB_INV8.I FULL_COUNTER.O.8 DC 0
V507 FULL_COUNTER.O.8 FULL_COUNTER.COUNT_SUB_DFF8.Q DC 0
V508 FULL_COUNTER.COUNT_SUB_DFF8.RSTb FULL_COUNTER.RSTb DC 0
V509 FULL_COUNTER.COUNT_SUB_DFF8.D FULL_COUNTER.D.8 DC 0
V510 FULL_COUNTER.COUNT_SUB_DFF8.CLK FULL_COUNTER.O.7 DC 0
V511 FULL_COUNTER.D.9 FULL_COUNTER.COUNT_SUB_INV9.O DC 0
V512 FULL_COUNTER.COUNT_SUB_INV9.I FULL_COUNTER.O.9 DC 0
V513 FULL_COUNTER.O.9 FULL_COUNTER.COUNT_SUB_DFF9.Q DC 0
V514 FULL_COUNTER.COUNT_SUB_DFF9.RSTb FULL_COUNTER.RSTb DC 0
V515 FULL_COUNTER.COUNT_SUB_DFF9.D FULL_COUNTER.D.9 DC 0
V516 FULL_COUNTER.COUNT_SUB_DFF9.CLK FULL_COUNTER.O.8 DC 0
V517 FULL_COUNTER.D.10 FULL_COUNTER.COUNT_SUB_INV10.O DC 0
V518 FULL_COUNTER.COUNT_SUB_INV10.I FULL_COUNTER.O.10 DC 0
V519 FULL_COUNTER.O.10 FULL_COUNTER.COUNT_SUB_DFF10.Q DC 0
V520 FULL_COUNTER.COUNT_SUB_DFF10.RSTb FULL_COUNTER.RSTb DC 0
V521 FULL_COUNTER.COUNT_SUB_DFF10.D FULL_COUNTER.D.10 DC 0
V522 FULL_COUNTER.COUNT_SUB_DFF10.CLK FULL_COUNTER.O.9 DC 0
V523 FULL_COUNTER.D.11 FULL_COUNTER.COUNT_SUB_INV11.O DC 0
V524 FULL_COUNTER.COUNT_SUB_INV11.I FULL_COUNTER.O.11 DC 0
V525 FULL_COUNTER.O.11 FULL_COUNTER.COUNT_SUB_DFF11.Q DC 0
V526 FULL_COUNTER.COUNT_SUB_DFF11.RSTb FULL_COUNTER.RSTb DC 0
V527 FULL_COUNTER.COUNT_SUB_DFF11.D FULL_COUNTER.D.11 DC 0
V528 FULL_COUNTER.COUNT_SUB_DFF11.CLK FULL_COUNTER.O.10 DC 0
V529 FULL_COUNTER.D.12 FULL_COUNTER.COUNT_SUB_INV12.O DC 0
V530 FULL_COUNTER.COUNT_SUB_INV12.I FULL_COUNTER.O.12 DC 0
V531 FULL_COUNTER.O.12 FULL_COUNTER.COUNT_SUB_DFF12.Q DC 0
V532 FULL_COUNTER.COUNT_SUB_DFF12.RSTb FULL_COUNTER.RSTb DC 0
V533 FULL_COUNTER.COUNT_SUB_DFF12.D FULL_COUNTER.D.12 DC 0
V534 FULL_COUNTER.COUNT_SUB_DFF12.CLK FULL_COUNTER.O.11 DC 0
V535 FULL_COUNTER.D.13 FULL_COUNTER.COUNT_SUB_INV13.O DC 0
V536 FULL_COUNTER.COUNT_SUB_INV13.I FULL_COUNTER.O.13 DC 0
V537 FULL_COUNTER.O.13 FULL_COUNTER.COUNT_SUB_DFF13.Q DC 0
V538 FULL_COUNTER.COUNT_SUB_DFF13.RSTb FULL_COUNTER.RSTb DC 0
V539 FULL_COUNTER.COUNT_SUB_DFF13.D FULL_COUNTER.D.13 DC 0
V540 FULL_COUNTER.COUNT_SUB_DFF13.CLK FULL_COUNTER.O.12 DC 0
V541 FULL_COUNTER.D.14 FULL_COUNTER.COUNT_SUB_INV14.O DC 0
V542 FULL_COUNTER.COUNT_SUB_INV14.I FULL_COUNTER.O.14 DC 0
V543 FULL_COUNTER.O.14 FULL_COUNTER.COUNT_SUB_DFF14.Q DC 0
V544 FULL_COUNTER.COUNT_SUB_DFF14.RSTb FULL_COUNTER.RSTb DC 0
V545 FULL_COUNTER.COUNT_SUB_DFF14.D FULL_COUNTER.D.14 DC 0
V546 FULL_COUNTER.COUNT_SUB_DFF14.CLK FULL_COUNTER.O.13 DC 0
V547 FULL_COUNTER.D.15 FULL_COUNTER.COUNT_SUB_INV15.O DC 0
V548 FULL_COUNTER.COUNT_SUB_INV15.I FULL_COUNTER.O.15 DC 0
V549 FULL_COUNTER.O.15 FULL_COUNTER.COUNT_SUB_DFF15.Q DC 0
V550 FULL_COUNTER.COUNT_SUB_DFF15.RSTb FULL_COUNTER.RSTb DC 0
V551 FULL_COUNTER.COUNT_SUB_DFF15.D FULL_COUNTER.D.15 DC 0
V552 FULL_COUNTER.COUNT_SUB_DFF15.CLK FULL_COUNTER.O.14 DC 0
V553 FULL_COUNTER.D.16 FULL_COUNTER.COUNT_SUB_INV16.O DC 0
V554 FULL_COUNTER.COUNT_SUB_INV16.I FULL_COUNTER.O.16 DC 0
V555 FULL_COUNTER.O.16 FULL_COUNTER.COUNT_SUB_DFF16.Q DC 0
V556 FULL_COUNTER.COUNT_SUB_DFF16.RSTb FULL_COUNTER.RSTb DC 0
V557 FULL_COUNTER.COUNT_SUB_DFF16.D FULL_COUNTER.D.16 DC 0
V558 FULL_COUNTER.COUNT_SUB_DFF16.CLK FULL_COUNTER.O.15 DC 0
V559 FULL_COUNTER.D.17 FULL_COUNTER.COUNT_SUB_INV17.O DC 0
V560 FULL_COUNTER.COUNT_SUB_INV17.I FULL_COUNTER.O.17 DC 0
V561 FULL_COUNTER.O.17 FULL_COUNTER.COUNT_SUB_DFF17.Q DC 0
V562 FULL_COUNTER.COUNT_SUB_DFF17.RSTb FULL_COUNTER.RSTb DC 0
V563 FULL_COUNTER.COUNT_SUB_DFF17.D FULL_COUNTER.D.17 DC 0
V564 FULL_COUNTER.COUNT_SUB_DFF17.CLK FULL_COUNTER.O.16 DC 0
V565 FULL_COUNTER.D.18 FULL_COUNTER.COUNT_SUB_INV18.O DC 0
V566 FULL_COUNTER.COUNT_SUB_INV18.I FULL_COUNTER.O.18 DC 0
V567 FULL_COUNTER.O.18 FULL_COUNTER.COUNT_SUB_DFF18.Q DC 0
V568 FULL_COUNTER.COUNT_SUB_DFF18.RSTb FULL_COUNTER.RSTb DC 0
V569 FULL_COUNTER.COUNT_SUB_DFF18.D FULL_COUNTER.D.18 DC 0
V570 FULL_COUNTER.COUNT_SUB_DFF18.CLK FULL_COUNTER.O.17 DC 0
V571 RISING_COUNTER.D.15 RISING_COUNTER.COUNT_SUB_INV15.O DC 0
V572 RISING_COUNTER.COUNT_SUB_INV15.I RISING_COUNTER.O.15 DC 0
V573 RISING_COUNTER.O.15 RISING_COUNTER.COUNT_SUB_DFF15.Q DC 0
V574 RISING_COUNTER.COUNT_SUB_DFF15.RSTb RISING_COUNTER.RSTb DC 0
V575 RISING_COUNTER.COUNT_SUB_DFF15.D RISING_COUNTER.D.15 DC 0
V576 RISING_COUNTER.COUNT_SUB_DFF15.CLK RISING_COUNTER.O.14 DC 0
V577 FULL_COUNTER.D.19 FULL_COUNTER.COUNT_SUB_INV19.O DC 0
V578 FULL_COUNTER.COUNT_SUB_INV19.I FULL_COUNTER.O.19 DC 0
V579 FULL_COUNTER.O.19 FULL_COUNTER.COUNT_SUB_DFF19.Q DC 0
V580 FULL_COUNTER.COUNT_SUB_DFF19.RSTb FULL_COUNTER.RSTb DC 0
V581 FULL_COUNTER.COUNT_SUB_DFF19.D FULL_COUNTER.D.19 DC 0
V582 FULL_COUNTER.COUNT_SUB_DFF19.CLK FULL_COUNTER.O.18 DC 0

.ends
