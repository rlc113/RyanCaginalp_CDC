* SPICE3 file created from SLC.ext - technology: sky130A

* .option scale=10n

.subckt SLC VGND VPB VNB INB IN VPWR VOUT
X0 VGND IN a_264_22# VNB sky130_fd_pr__nfet_01v8_lvt ad=135 pd=15.4 as=72.5 ps=7.9 w=5e+07 l=1.5e+07 M=10
X1 a_919_243# INB VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=72.5 pd=7.9 as=72.5 ps=7.9 w=5e+07 l=1.5e+07 M=10
X2 a_438_293# a_264_22# a_264_22# VPB sky130_fd_pr__pfet_01v8_hvt ad=522 pd=65 as=972 ps=126 w=3.6e+07 l=1.5e+07
X3 VPWR a_438_293# VOUT VPB sky130_fd_pr__pfet_01v8_hvt ad=762 pd=80.5 as=362 ps=39.5 w=5e+07 l=1.5e+07 M=2
X4 VGND a_264_22# VOUT VNB sky130_fd_pr__nfet_01v8 ad=1.75k pd=184 as=1.75k ps=184 w=6.5e+07 l=1.5e+07
X5 a_1235_416# a_264_22# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=522 pd=65 as=972 ps=126 w=3.6e+07 l=1.5e+07
X6 VPWR a_919_243# a_438_293# VPB sky130_fd_pr__pfet_01v8_hvt ad=972 pd=126 as=522 ps=65 w=3.6e+07 l=1.5e+07
X7 a_919_243# a_919_243# a_1235_416# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.12k pd=134 as=522 ps=65 w=3.6e+07 l=1.5e+07
.ends
