* NGSPICE file created from CDC.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_16 VNB VPB VGND VPWR Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 Y VPB 0.0305f
C1 VPWR A 0.28f
C2 Y VGND 1.06f
C3 VPWR VPB 0.159f
C4 VPB A 0.526f
C5 VGND VPWR 0.161f
C6 VGND A 0.266f
C7 Y VPWR 1.47f
C8 Y A 1.43f
C9 VGND VPB 0.0132f
C10 VGND VNB 0.865f
C11 Y VNB 0.0551f
C12 VPWR VNB 0.737f
C13 A VNB 1.55f
C14 VPB VNB 1.49f
.ends

.subckt sky130_fd_sc_hd__nand2_8 VNB VPB VGND VPWR A Y B a_27_47#
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VPWR Y 1.49f
C1 B VPB 0.248f
C2 B VGND 0.108f
C3 VPB VGND 0.0101f
C4 Y a_27_47# 0.337f
C5 A Y 0.644f
C6 VPWR a_27_47# 0.0392f
C7 A VPWR 0.129f
C8 Y B 0.413f
C9 A a_27_47# 0.0695f
C10 Y VPB 0.0366f
C11 Y VGND 0.0559f
C12 VPWR B 0.118f
C13 VPWR VPB 0.157f
C14 VPWR VGND 0.149f
C15 B a_27_47# 0.369f
C16 A B 0.051f
C17 VPB a_27_47# 0.00278f
C18 VGND a_27_47# 0.947f
C19 A VPB 0.247f
C20 A VGND 0.0645f
C21 VGND VNB 0.797f
C22 Y VNB 0.0446f
C23 VPWR VNB 0.753f
C24 A VNB 0.746f
C25 B VNB 0.758f
C26 VPB VNB 1.49f
C27 a_27_47# VNB 0.083f
.ends

.subckt transmission_gate G VPWR VGND O GN
X0 O G VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.226 pd=1.92 as=0.226 ps=1.92 w=0.55 l=0.15
X1 O GN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.226 pd=1.92 as=0.226 ps=1.92 w=0.55 l=0.15
C0 GN VPWR 0.26f
C1 O G 0.0806f
C2 G GN 0.0779f
C3 G VPWR 0.0769f
C4 O GN 0.0362f
C5 O VPWR 0.154f
C6 G VGND 0.21f
C7 O VGND 0.13f
C8 GN VGND 0.0906f
C9 VPWR VGND 1.26f
.ends

.subckt sky130_fd_sc_hd__decap_4 VNB VPB VGND VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VGND VPWR 0.546f
C1 VPWR VPB 0.0787f
C2 VGND VPB 0.116f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__dfbbn_1 VNB VPB VGND VPWR Q Q_N RESET_B SET_B D CLK_N a_2136_47#
+ a_791_47# a_647_21# a_891_329# a_1363_47# a_557_413# a_941_21# a_1415_315# a_473_413#
+ a_193_47# a_381_47# a_1112_329# a_1555_47# a_581_47# a_1340_413# a_1159_47# a_1256_413#
+ a_1672_329# a_27_47#
X0 a_791_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1 a_1555_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2 VPWR RESET_B a_941_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X3 a_1415_315# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X4 a_791_47# a_941_21# a_647_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VGND a_1415_315# a_1363_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X6 a_1340_413# a_27_47# a_1256_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_473_413# a_193_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X10 a_1555_47# a_941_21# a_1415_315# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VPWR a_1415_315# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_1256_413# a_193_47# a_1112_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X13 a_581_47# a_27_47# a_473_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X14 a_647_21# a_473_413# a_791_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X15 a_647_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X16 VPWR a_941_21# a_891_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X17 a_557_413# a_193_47# a_473_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X20 a_473_413# a_27_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X21 a_891_329# a_473_413# a_647_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X22 Q_N a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X23 VGND RESET_B a_941_21# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X24 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X25 VPWR a_647_21# a_557_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X26 a_1112_329# a_647_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X27 VGND a_647_21# a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X28 VGND a_1415_315# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 VPWR a_941_21# a_1672_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X31 VPWR a_1415_315# a_1340_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X32 a_1363_47# a_193_47# a_1256_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X33 Q_N a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X35 a_1159_47# a_647_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X36 a_1672_329# a_1256_413# a_1415_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X37 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X38 a_1256_413# a_27_47# a_1159_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X39 a_1415_315# a_1256_413# a_1555_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
C0 a_647_21# a_1159_47# 9.75e-19
C1 a_647_21# VGND 0.053f
C2 a_193_47# a_557_413# 0.0018f
C3 a_27_47# a_891_329# 2.46e-19
C4 a_791_47# a_1159_47# 3.34e-19
C5 a_381_47# VGND 0.0775f
C6 a_791_47# VGND 0.164f
C7 a_27_47# D 0.11f
C8 a_2136_47# Q 0.0721f
C9 a_1555_47# SET_B 0.0131f
C10 a_2136_47# VPWR 0.139f
C11 a_193_47# a_1159_47# 2.14e-20
C12 VPB CLK_N 0.0706f
C13 a_1159_47# a_1256_413# 0.00386f
C14 a_941_21# VPB 0.142f
C15 a_193_47# VGND 0.0661f
C16 VGND Q_N 0.0862f
C17 a_1256_413# VGND 0.127f
C18 a_941_21# a_1415_315# 0.267f
C19 a_647_21# RESET_B 6.51e-21
C20 a_381_47# RESET_B 3.34e-21
C21 a_27_47# SET_B 0.309f
C22 a_381_47# a_647_21# 8.07e-20
C23 a_941_21# a_1112_329# 0.00652f
C24 a_2136_47# VGND 0.114f
C25 a_647_21# a_791_47# 0.0697f
C26 a_1555_47# VPWR 1.3e-19
C27 a_1363_47# SET_B 7.87e-19
C28 VPB D 0.0817f
C29 a_941_21# CLK_N 5.45e-20
C30 a_193_47# RESET_B 6.8e-20
C31 RESET_B Q_N 0.0017f
C32 a_1256_413# RESET_B 4.43e-20
C33 a_1340_413# VPWR 0.00281f
C34 a_473_413# a_27_47# 0.159f
C35 a_647_21# a_193_47# 0.117f
C36 a_647_21# a_1256_413# 0.00189f
C37 a_381_47# a_193_47# 0.189f
C38 a_193_47# a_791_47# 6.04e-20
C39 a_27_47# a_581_47# 0.00206f
C40 a_27_47# Q 2.71e-20
C41 a_791_47# a_1256_413# 0.00316f
C42 a_27_47# VPWR 0.146f
C43 a_941_21# a_891_329# 1.21e-20
C44 a_193_47# a_1672_329# 7.17e-20
C45 a_1555_47# VGND 0.157f
C46 a_2136_47# RESET_B 4.99e-19
C47 a_1672_329# Q_N 2.1e-20
C48 VPB SET_B 0.147f
C49 a_941_21# D 1.12e-19
C50 a_193_47# Q_N 1.07e-19
C51 a_27_47# a_557_413# 4.45e-20
C52 a_193_47# a_1256_413# 0.0334f
C53 a_1256_413# Q_N 1e-20
C54 a_1415_315# SET_B 0.141f
C55 a_27_47# a_1159_47# 0.00272f
C56 a_473_413# VPB 0.0627f
C57 a_27_47# VGND 0.292f
C58 a_473_413# a_1415_315# 4.59e-22
C59 a_193_47# a_2136_47# 1.03e-19
C60 a_1363_47# VGND 0.00192f
C61 a_1555_47# RESET_B 3.78e-20
C62 a_2136_47# Q_N 0.175f
C63 Q VPB 0.0123f
C64 VPB VPWR 0.255f
C65 a_941_21# SET_B 0.096f
C66 a_1415_315# Q 0.00311f
C67 a_1415_315# VPWR 0.315f
C68 a_27_47# RESET_B 2.12e-19
C69 a_473_413# a_941_21# 0.0633f
C70 a_1112_329# VPWR 0.0164f
C71 a_1555_47# a_1256_413# 0.0256f
C72 a_647_21# a_27_47# 0.15f
C73 a_941_21# Q 1.7e-19
C74 VPB VGND 0.0151f
C75 CLK_N VPWR 0.0196f
C76 a_941_21# VPWR 0.197f
C77 a_381_47# a_27_47# 0.0456f
C78 a_1415_315# VGND 0.0797f
C79 a_27_47# a_791_47# 0.00134f
C80 a_1340_413# a_1256_413# 0.00857f
C81 a_1363_47# a_791_47# 2.46e-21
C82 a_473_413# D 1.43e-19
C83 a_27_47# a_193_47# 0.798f
C84 a_27_47# Q_N 4.78e-20
C85 a_27_47# a_1256_413# 0.14f
C86 a_891_329# VPWR 0.00984f
C87 a_1112_329# VGND 3.84e-19
C88 a_1363_47# a_1256_413# 0.00707f
C89 a_941_21# a_1159_47# 3.73e-19
C90 CLK_N VGND 0.0196f
C91 D VPWR 0.0153f
C92 VPB RESET_B 0.0476f
C93 a_941_21# VGND 0.134f
C94 a_1415_315# RESET_B 0.0851f
C95 a_647_21# VPB 0.141f
C96 a_381_47# VPB 0.0197f
C97 a_27_47# a_2136_47# 1.76e-19
C98 a_473_413# SET_B 0.14f
C99 Q SET_B 1.24e-19
C100 a_193_47# VPB 0.198f
C101 SET_B VPWR 0.0255f
C102 D VGND 0.0134f
C103 VPB Q_N 0.0102f
C104 a_1256_413# VPB 0.0597f
C105 a_1415_315# a_1672_329# 0.00869f
C106 a_941_21# RESET_B 0.105f
C107 a_647_21# a_1112_329# 9.46e-19
C108 a_1415_315# a_193_47# 0.0494f
C109 a_1415_315# Q_N 0.121f
C110 a_1415_315# a_1256_413# 0.207f
C111 a_941_21# a_647_21# 0.199f
C112 a_941_21# a_381_47# 3.79e-20
C113 a_473_413# a_581_47# 0.00807f
C114 a_941_21# a_791_47# 0.00926f
C115 a_473_413# VPWR 0.108f
C116 a_1555_47# a_1363_47# 4.19e-20
C117 a_27_47# a_1340_413# 2.13e-19
C118 a_193_47# a_1112_329# 0.00907f
C119 a_2136_47# VPB 0.0467f
C120 a_1112_329# a_1256_413# 0.00412f
C121 a_941_21# a_1672_329# 0.0016f
C122 a_1159_47# SET_B 0.00459f
C123 Q VPWR 0.0992f
C124 a_193_47# CLK_N 7.87e-19
C125 SET_B VGND 0.311f
C126 a_1415_315# a_2136_47# 0.0967f
C127 a_941_21# a_193_47# 0.126f
C128 a_941_21# Q_N 0.0054f
C129 a_941_21# a_1256_413# 0.13f
C130 a_473_413# a_557_413# 0.00972f
C131 a_647_21# a_891_329# 0.0104f
C132 a_557_413# VPWR 0.0042f
C133 a_381_47# D 0.148f
C134 a_473_413# VGND 0.147f
C135 a_193_47# a_891_329# 0.00276f
C136 a_1555_47# VPB 8.96e-20
C137 a_941_21# a_2136_47# 5.84e-19
C138 a_1159_47# VPWR 6.2e-19
C139 a_581_47# VGND 0.0017f
C140 Q VGND 0.0643f
C141 a_193_47# D 0.0986f
C142 VPWR VGND 0.0801f
C143 SET_B RESET_B 0.00229f
C144 a_1415_315# a_1555_47# 0.0383f
C145 a_647_21# SET_B 0.175f
C146 a_791_47# SET_B 0.03f
C147 a_27_47# VPB 0.224f
C148 a_473_413# RESET_B 7.48e-21
C149 a_1415_315# a_27_47# 0.0321f
C150 a_941_21# a_1555_47# 0.0526f
C151 a_1159_47# VGND 0.0108f
C152 Q RESET_B 6.25e-20
C153 a_473_413# a_647_21# 0.206f
C154 a_193_47# SET_B 0.0123f
C155 VPWR RESET_B 0.0099f
C156 SET_B Q_N 3.72e-19
C157 a_1256_413# SET_B 0.177f
C158 a_473_413# a_381_47# 0.0369f
C159 a_941_21# a_1340_413# 9.41e-19
C160 a_473_413# a_791_47# 0.025f
C161 a_647_21# VPWR 0.16f
C162 a_381_47# a_581_47# 3.81e-19
C163 a_27_47# a_1112_329# 1.09e-19
C164 a_381_47# VPWR 0.0894f
C165 a_27_47# CLK_N 0.212f
C166 a_941_21# a_27_47# 0.14f
C167 a_473_413# a_193_47# 0.15f
C168 a_647_21# a_557_413# 6.69e-20
C169 a_2136_47# SET_B 3.22e-19
C170 a_1672_329# VPWR 0.00438f
C171 a_941_21# a_1363_47# 1.96e-20
C172 a_381_47# a_557_413# 8.99e-19
C173 a_193_47# Q 5.52e-20
C174 a_193_47# VPWR 0.443f
C175 VPWR Q_N 0.0614f
C176 VGND RESET_B 0.0282f
C177 a_1256_413# VPWR 0.12f
C178 a_1415_315# VPB 0.242f
C179 Q VNB 0.0945f
C180 Q_N VNB 0.0135f
C181 RESET_B VNB 0.133f
C182 VGND VNB 1.3f
C183 VPWR VNB 1.05f
C184 SET_B VNB 0.264f
C185 D VNB 0.125f
C186 CLK_N VNB 0.197f
C187 VPB VNB 2.38f
C188 a_1555_47# VNB 0.00871f
C189 a_2136_47# VNB 0.133f
C190 a_791_47# VNB 0.0125f
C191 a_381_47# VNB 0.0218f
C192 a_1256_413# VNB 0.12f
C193 a_1415_315# VNB 0.394f
C194 a_941_21# VNB 0.245f
C195 a_473_413# VNB 0.119f
C196 a_647_21# VNB 0.24f
C197 a_193_47# VNB 0.27f
C198 a_27_47# VNB 0.492f
.ends

.subckt sky130_fd_sc_hd__inv_1 VNB VPB VGND VPWR A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
C0 A Y 0.0476f
C1 VPWR Y 0.128f
C2 VGND VPB 0.00948f
C3 VGND A 0.04f
C4 VPB A 0.0451f
C5 VGND VPWR 0.0338f
C6 VPB VPWR 0.0545f
C7 VGND Y 0.0998f
C8 VPB Y 0.0177f
C9 A VPWR 0.037f
C10 VGND VNB 0.251f
C11 Y VNB 0.0961f
C12 VPWR VNB 0.219f
C13 A VNB 0.167f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__inv_8 VNB VPB VGND VPWR Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 A Y 0.829f
C1 VPWR Y 0.78f
C2 VGND VPB 0.00793f
C3 VGND A 0.117f
C4 VPB A 0.254f
C5 VGND VPWR 0.0854f
C6 VPB VPWR 0.1f
C7 VGND Y 0.574f
C8 VPB Y 0.0348f
C9 A VPWR 0.128f
C10 VGND VNB 0.51f
C11 Y VNB 0.127f
C12 VPWR VNB 0.45f
C13 A VNB 0.771f
C14 VPB VNB 0.871f
.ends

.subckt sky130_fd_sc_hd__nor2_1 VNB VPB VGND VPWR A B Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB A 0.0415f
C1 VPWR a_109_297# 0.00638f
C2 B A 0.0584f
C3 VGND VPWR 0.0314f
C4 Y VPWR 0.0995f
C5 VPWR VPB 0.0449f
C6 VGND a_109_297# 0.00128f
C7 Y a_109_297# 0.0113f
C8 VPWR B 0.0148f
C9 VPWR A 0.0528f
C10 VGND Y 0.154f
C11 VGND VPB 0.00456f
C12 Y VPB 0.0139f
C13 VGND B 0.0451f
C14 Y B 0.0877f
C15 VGND A 0.0486f
C16 Y A 0.0471f
C17 VPB B 0.0367f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__inv_4 VNB VPB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VGND VPWR 0.0501f
C1 VPB VPWR 0.0654f
C2 A VGND 0.0819f
C3 A VPB 0.142f
C4 VGND VPB 0.00667f
C5 Y VPWR 0.362f
C6 A Y 0.36f
C7 VGND Y 0.263f
C8 Y VPB 0.0159f
C9 A VPWR 0.0982f
C10 VGND VNB 0.327f
C11 Y VNB 0.0849f
C12 VPWR VNB 0.296f
C13 A VNB 0.452f
C14 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__inv_2 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 VGND VPWR 0.0423f
C1 VPB VPWR 0.0521f
C2 A VGND 0.0638f
C3 A VPB 0.0742f
C4 VGND VPB 0.00649f
C5 Y VPWR 0.209f
C6 A Y 0.0894f
C7 VGND Y 0.155f
C8 Y VPB 0.0061f
C9 A VPWR 0.0631f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__conb_1 VNB VPB VGND VPWR LO HI
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
C0 VPB VGND 0.00479f
C1 VPWR HI 0.0726f
C2 VPWR LO 0.241f
C3 VPWR VGND 0.0317f
C4 VPB VPWR 0.158f
C5 HI LO 0.0683f
C6 HI VGND 0.207f
C7 VPB HI 0.00473f
C8 LO VGND 0.0605f
C9 VPB LO 0.134f
C10 VGND VNB 0.406f
C11 LO VNB 0.166f
C12 HI VNB 0.25f
C13 VPWR VNB 0.297f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nand3_1 VNB VPB VGND VPWR A B Y C a_193_47# a_109_47#
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y a_193_47# 0.0117f
C1 Y A 0.0909f
C2 VPB C 0.0373f
C3 VGND VPB 0.00519f
C4 a_109_47# VGND 9.04e-19
C5 VGND C 0.0415f
C6 VPWR a_193_47# 5.03e-19
C7 B a_193_47# 0.00347f
C8 VPWR A 0.0186f
C9 VPWR Y 0.317f
C10 B A 0.0823f
C11 Y B 0.149f
C12 A VPB 0.0368f
C13 VGND a_193_47# 0.00142f
C14 Y VPB 0.0166f
C15 VPWR B 0.017f
C16 A VGND 0.01f
C17 Y a_109_47# 0.0108f
C18 Y C 0.0724f
C19 Y VGND 0.181f
C20 VPWR VPB 0.0506f
C21 B VPB 0.0268f
C22 VPWR a_109_47# 2.94e-19
C23 VPWR C 0.0414f
C24 VPWR VGND 0.0416f
C25 a_109_47# B 4.42e-19
C26 B C 0.051f
C27 B VGND 0.0116f
C28 VGND VNB 0.263f
C29 Y VNB 0.0816f
C30 VPWR VNB 0.247f
C31 A VNB 0.143f
C32 B VNB 0.0976f
C33 C VNB 0.157f
C34 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__nand2_1 VNB VPB VGND VPWR A Y B a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 VGND VPWR 0.0322f
C1 VPWR Y 0.211f
C2 B VPWR 0.0478f
C3 A VGND 0.00949f
C4 A Y 0.0855f
C5 A B 0.051f
C6 VGND Y 0.139f
C7 VGND B 0.0544f
C8 B Y 0.0481f
C9 VPB VPWR 0.0509f
C10 VPB A 0.0379f
C11 VPB VGND 0.0044f
C12 VPB Y 0.00618f
C13 VPB B 0.0391f
C14 a_113_47# VPWR 1.78e-19
C15 VGND a_113_47# 0.0019f
C16 A VPWR 0.0444f
C17 a_113_47# Y 0.00937f
C18 VGND VNB 0.232f
C19 Y VNB 0.0557f
C20 VPWR VNB 0.245f
C21 A VNB 0.143f
C22 B VNB 0.146f
C23 VPB VNB 0.339f
.ends

.subckt CDC Reset CLOCK_GEN.SR_Op.Q V_GND V_LOW V_HIGH V_SENSE RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_DFF19.Q
Xsky130_fd_sc_hd__inv_16_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_16_3/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand3_1_2/Y CLOCK_GEN.SR_Op.Q
+ sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_31 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_20 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_75 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_53 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_42 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_64 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_90 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_6 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_10/HI
+ sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__dfbbn_1_6/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# sky130_fd_sc_hd__dfbbn_1_6/a_557_413# sky130_fd_sc_hd__dfbbn_1_6/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__dfbbn_1_6/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_581_47# sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# sky130_fd_sc_hd__dfbbn_1_6/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# sky130_fd_sc_hd__dfbbn_1_6/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_4 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_4/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_15 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF17.Q
+ sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_48 V_GND V_LOW V_GND V_LOW Reset sky130_fd_sc_hd__inv_1_48/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_37 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_26 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_59 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__inv_1_59/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_8_0/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_64/A
+ sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_32 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_10 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_21 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_43 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_65 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_54 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_76 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_91 V_GND sky130_fd_sc_hd__fill_8_848/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 V_GND sky130_fd_sc_hd__fill_8_949/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_7 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_5/HI
+ sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_7/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# sky130_fd_sc_hd__dfbbn_1_7/a_557_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# sky130_fd_sc_hd__dfbbn_1_7/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_581_47# sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# sky130_fd_sc_hd__dfbbn_1_7/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# sky130_fd_sc_hd__dfbbn_1_7/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_5 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_5/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_16 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF19.Q
+ sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_27 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_49 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_38 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__inv_1_38/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_16_5/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__nand2_8_4/Y
+ CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_22 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_11 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_44 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_33 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_55 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_66 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_77 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_70 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 V_GND sky130_fd_sc_hd__fill_8_949/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_92 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_8 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_8/HI
+ sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__dfbbn_1_8/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_8/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# sky130_fd_sc_hd__dfbbn_1_8/a_557_413# sky130_fd_sc_hd__dfbbn_1_8/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_8/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# sky130_fd_sc_hd__dfbbn_1_8/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_581_47# sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# sky130_fd_sc_hd__dfbbn_1_8/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# sky130_fd_sc_hd__dfbbn_1_8/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_6 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_6/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_17 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_67/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_39 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_28 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_6/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_56/Y sky130_fd_sc_hd__inv_1_53/A
+ sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__inv_8_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_8_0/A
+ sky130_fd_sc_hd__inv_8
Xtransmission_gate_23 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_12 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_45 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_34 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_56 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_67 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_78 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_60 V_GND sky130_fd_sc_hd__fill_8_848/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 V_GND sky130_fd_sc_hd__fill_8_927/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 V_GND sky130_fd_sc_hd__fill_8_951/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_9 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_6/HI
+ sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__dfbbn_1_9/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# sky130_fd_sc_hd__dfbbn_1_9/a_557_413# sky130_fd_sc_hd__dfbbn_1_9/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# sky130_fd_sc_hd__dfbbn_1_9/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_581_47# sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# sky130_fd_sc_hd__dfbbn_1_9/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# sky130_fd_sc_hd__dfbbn_1_9/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_7 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_7/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_18 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_18/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_29 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_52/A
+ sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_13 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_46 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_24 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_57 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_35 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_79 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_68 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_50 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 V_GND sky130_fd_sc_hd__fill_8_854/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_72 V_GND sky130_fd_sc_hd__fill_8_958/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 V_GND sky130_fd_sc_hd__fill_8_951/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_8 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_8/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_19 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_19/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_50 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_50/Y
+ sky130_fd_sc_hd__inv_16_50/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_8/Y sky130_fd_sc_hd__inv_16_8/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_65/A
+ sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_14 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_47 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_36 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_25 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_58 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_69 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_51 V_GND sky130_fd_sc_hd__fill_8_858/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_40 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_62 V_GND sky130_fd_sc_hd__fill_8_858/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_73 V_GND sky130_fd_sc_hd__fill_8_927/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 V_GND sky130_fd_sc_hd__fill_8_949/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_95 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_9 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_9/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor2_1_0 V_GND V_LOW V_GND V_LOW Reset CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__inv_16_40 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_40/Y Reset
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_51 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_51/Y
+ sky130_fd_sc_hd__inv_16_51/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_9/Y sky130_fd_sc_hd__inv_16_9/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_47/A
+ sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_37 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_26 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_15 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_48 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_59 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_30 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_52 V_GND sky130_fd_sc_hd__fill_8_852/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_63 V_GND sky130_fd_sc_hd__fill_8_858/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 V_GND sky130_fd_sc_hd__fill_8_951/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_96 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_30 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_16_31/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_52 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_46/A
+ sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_41 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_41/Y Reset
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__nand2_8_9/Y
+ sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_38 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_16 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_27 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_49 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_20 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_53 V_GND sky130_fd_sc_hd__fill_8_848/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 V_GND sky130_fd_sc_hd__fill_8_927/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 V_GND sky130_fd_sc_hd__fill_8_927/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 V_GND sky130_fd_sc_hd__fill_8_949/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_97 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_31 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_1_67/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_20 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_16_20/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_53 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16_4/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_42 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_42/Y Reset
+ sky130_fd_sc_hd__inv_16
Xtransmission_gate_28 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_17 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_39 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_10 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 V_GND sky130_fd_sc_hd__fill_8_854/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_76 V_GND sky130_fd_sc_hd__fill_8_932/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 V_GND sky130_fd_sc_hd__fill_8_958/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_170 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_10 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_8/A sky130_fd_sc_hd__inv_16_28/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_21 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_22/A sky130_fd_sc_hd__inv_16_27/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_54 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__inv_16_6/A
+ sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_32 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_32/Y sky130_fd_sc_hd__inv_16_32/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_43 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_24/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_50 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_30/HI
+ sky130_fd_sc_hd__inv_1_38/Y RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__dfbbn_1_50/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_50/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# sky130_fd_sc_hd__dfbbn_1_50/a_557_413# sky130_fd_sc_hd__dfbbn_1_50/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_50/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# sky130_fd_sc_hd__dfbbn_1_50/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_581_47# sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# sky130_fd_sc_hd__dfbbn_1_50/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_50/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xtransmission_gate_18 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_29 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_11 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 V_GND sky130_fd_sc_hd__fill_8_852/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_77 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_88 V_GND sky130_fd_sc_hd__fill_8_958/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_99 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_160 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_171 V_GND sky130_fd_sc_hd__fill_4_320/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_4_0 V_GND V_LOW V_LOW V_GND sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_4_0/A
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_16_11 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_6/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_22 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_22/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_55 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_55/Y
+ sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_44 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_44/Y
+ sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_33 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_9/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_40 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_44/HI
+ sky130_fd_sc_hd__inv_1_60/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_40/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_40/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# sky130_fd_sc_hd__dfbbn_1_40/a_557_413# sky130_fd_sc_hd__dfbbn_1_40/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_40/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# sky130_fd_sc_hd__dfbbn_1_40/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_581_47# sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# sky130_fd_sc_hd__dfbbn_1_40/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_40/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_51 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_48/HI
+ sky130_fd_sc_hd__inv_1_59/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_51/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__dfbbn_1_51/a_557_413# sky130_fd_sc_hd__dfbbn_1_51/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_51/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__dfbbn_1_51/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_581_47# sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# sky130_fd_sc_hd__dfbbn_1_51/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_51/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xtransmission_gate_19 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_12 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 V_GND sky130_fd_sc_hd__fill_8_854/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_45 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_78 V_GND sky130_fd_sc_hd__fill_8_932/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_89 V_GND sky130_fd_sc_hd__fill_8_848/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 V_GND sky130_fd_sc_hd__fill_8_958/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_150 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_161 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_172 V_GND sky130_fd_sc_hd__fill_4_320/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_12 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_15/A sky130_fd_sc_hd__inv_16_14/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_45 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_55/A
+ sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_34 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_49/A
+ sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_56 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__inv_16_6/A
+ sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_23 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_16_23/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_30 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_28/HI
+ sky130_fd_sc_hd__inv_1_40/Y RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_30/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__dfbbn_1_30/a_557_413# sky130_fd_sc_hd__dfbbn_1_30/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_581_47# sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# sky130_fd_sc_hd__dfbbn_1_30/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_41 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_47/HI
+ sky130_fd_sc_hd__inv_1_57/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_41/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_41/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# sky130_fd_sc_hd__dfbbn_1_41/a_557_413# sky130_fd_sc_hd__dfbbn_1_41/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_41/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# sky130_fd_sc_hd__dfbbn_1_41/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_581_47# sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# sky130_fd_sc_hd__dfbbn_1_41/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_41/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__decap_4_13 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 V_GND sky130_fd_sc_hd__fill_8_854/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_46 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_68 V_GND sky130_fd_sc_hd__fill_8_932/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_79 V_GND sky130_fd_sc_hd__fill_8_951/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_140 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_162 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_151 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_173 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_13 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_15/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_35 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_51/A
+ sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_46 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_52/A
+ sky130_fd_sc_hd__inv_16_55/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_24 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_24/Y sky130_fd_sc_hd__inv_16_26/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_20 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_18/HI
+ sky130_fd_sc_hd__inv_1_27/Y RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_20/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# sky130_fd_sc_hd__dfbbn_1_20/a_557_413# sky130_fd_sc_hd__dfbbn_1_20/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__dfbbn_1_20/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# sky130_fd_sc_hd__dfbbn_1_20/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_581_47# sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# sky130_fd_sc_hd__dfbbn_1_20/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_20/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_31 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_34/HI
+ sky130_fd_sc_hd__inv_1_35/Y RISING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_31/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_31/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__dfbbn_1_31/a_557_413# sky130_fd_sc_hd__dfbbn_1_31/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_31/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__dfbbn_1_31/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_581_47# sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# sky130_fd_sc_hd__dfbbn_1_31/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_31/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_42 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_49/HI
+ sky130_fd_sc_hd__inv_1_63/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__dfbbn_1_42/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__dfbbn_1_42/a_557_413# sky130_fd_sc_hd__dfbbn_1_42/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# sky130_fd_sc_hd__dfbbn_1_42/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_581_47# sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# sky130_fd_sc_hd__dfbbn_1_42/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_42/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__decap_4_14 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 V_GND sky130_fd_sc_hd__fill_8_858/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_36 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 V_GND sky130_fd_sc_hd__fill_8_932/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 V_GND sky130_fd_sc_hd__fill_8_852/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_141 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_130 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_163 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_152 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_47 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_47/Y
+ sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_36 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_44/A
+ sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_14 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_16/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_25 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_29/A sky130_fd_sc_hd__inv_16_7/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_2_0 V_GND V_LOW V_LOW V_GND sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_2_0/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfbbn_1_10 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF17.Q
+ sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_13/HI
+ sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__dfbbn_1_10/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_10/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# sky130_fd_sc_hd__dfbbn_1_10/a_557_413# sky130_fd_sc_hd__dfbbn_1_10/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_10/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# sky130_fd_sc_hd__dfbbn_1_10/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_581_47# sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# sky130_fd_sc_hd__dfbbn_1_10/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_10/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_32 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_29/HI
+ sky130_fd_sc_hd__inv_1_34/Y RISING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# sky130_fd_sc_hd__dfbbn_1_32/a_557_413# sky130_fd_sc_hd__dfbbn_1_32/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_32/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# sky130_fd_sc_hd__dfbbn_1_32/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_581_47# sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# sky130_fd_sc_hd__dfbbn_1_32/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_32/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_21 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_22/HI
+ sky130_fd_sc_hd__inv_1_29/Y FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__dfbbn_1_21/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_21/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# sky130_fd_sc_hd__dfbbn_1_21/a_557_413# sky130_fd_sc_hd__dfbbn_1_21/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_21/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__dfbbn_1_21/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_581_47# sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# sky130_fd_sc_hd__dfbbn_1_21/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_21/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_43 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_46/HI
+ sky130_fd_sc_hd__inv_1_62/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_43/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# sky130_fd_sc_hd__dfbbn_1_43/a_557_413# sky130_fd_sc_hd__dfbbn_1_43/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# sky130_fd_sc_hd__dfbbn_1_43/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_581_47# sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# sky130_fd_sc_hd__dfbbn_1_43/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__decap_4_15 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 V_GND sky130_fd_sc_hd__fill_8_852/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xtransmission_gate_0 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_120 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_131 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_142 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_164 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_153 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_37 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_48/A
+ sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_15 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_15/Y sky130_fd_sc_hd__inv_16_15/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_26 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_26/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_48 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_48/Y
+ sky130_fd_sc_hd__inv_16_48/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_11 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF18.Q
+ sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_14/HI
+ sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__dfbbn_1_11/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_11/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_581_47# sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# sky130_fd_sc_hd__dfbbn_1_11/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_11/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_33 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_27/HI
+ sky130_fd_sc_hd__inv_1_36/Y RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_33/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# sky130_fd_sc_hd__dfbbn_1_33/a_557_413# sky130_fd_sc_hd__dfbbn_1_33/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_581_47# sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# sky130_fd_sc_hd__dfbbn_1_33/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_22 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_26/HI
+ sky130_fd_sc_hd__inv_1_31/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__dfbbn_1_22/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_22/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# sky130_fd_sc_hd__dfbbn_1_22/a_557_413# sky130_fd_sc_hd__dfbbn_1_22/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_22/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__dfbbn_1_22/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_581_47# sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# sky130_fd_sc_hd__dfbbn_1_22/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_22/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_44 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_33/HI
+ sky130_fd_sc_hd__inv_1_39/Y RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# sky130_fd_sc_hd__dfbbn_1_44/a_557_413# sky130_fd_sc_hd__dfbbn_1_44/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# sky130_fd_sc_hd__dfbbn_1_44/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_581_47# sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# sky130_fd_sc_hd__dfbbn_1_44/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_50 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_50/LO
+ sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_16 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_38 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xtransmission_gate_1 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_121 V_GND sky130_fd_sc_hd__fill_4_188/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_132 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_110 V_GND sky130_fd_sc_hd__fill_4_182/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_143 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_165 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_154 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_38 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_45/A
+ sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_16 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_16/Y sky130_fd_sc_hd__inv_16_33/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_27 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_29/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_49 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_49/Y
+ sky130_fd_sc_hd__inv_16_49/A sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_12 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF19.Q
+ sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_11/HI
+ sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF18.Q sky130_fd_sc_hd__dfbbn_1_12/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# sky130_fd_sc_hd__dfbbn_1_12/a_557_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_581_47# sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# sky130_fd_sc_hd__dfbbn_1_12/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_23 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_50/HI
+ sky130_fd_sc_hd__inv_1_58/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__dfbbn_1_23/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# sky130_fd_sc_hd__dfbbn_1_23/a_557_413# sky130_fd_sc_hd__dfbbn_1_23/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# sky130_fd_sc_hd__dfbbn_1_23/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_34 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_51/HI
+ sky130_fd_sc_hd__inv_1_42/Y FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_34/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_34/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__dfbbn_1_34/a_557_413# sky130_fd_sc_hd__dfbbn_1_34/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_34/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# sky130_fd_sc_hd__dfbbn_1_34/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# sky130_fd_sc_hd__dfbbn_1_34/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_34/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_45 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_38/HI
+ sky130_fd_sc_hd__inv_1_49/Y RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_45/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# sky130_fd_sc_hd__dfbbn_1_45/a_557_413# sky130_fd_sc_hd__dfbbn_1_45/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# sky130_fd_sc_hd__dfbbn_1_45/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_581_47# sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# sky130_fd_sc_hd__dfbbn_1_45/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__dfbbn_1_45/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_40 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_40/LO
+ sky130_fd_sc_hd__conb_1_40/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_51 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_51/LO
+ sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_17 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xtransmission_gate_2 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_122 V_GND sky130_fd_sc_hd__fill_4_189/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_100 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_111 V_GND sky130_fd_sc_hd__fill_4_184/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_155 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_133 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_144 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_166 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_28 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_28/Y sky130_fd_sc_hd__inv_16_32/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_17 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_20/A sky130_fd_sc_hd__inv_16_24/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_39 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_16_50/A
+ sky130_fd_sc_hd__inv_16_51/Y sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_13 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF16.Q
+ sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_15/HI
+ sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_13/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# sky130_fd_sc_hd__dfbbn_1_13/a_557_413# sky130_fd_sc_hd__dfbbn_1_13/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_581_47# sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# sky130_fd_sc_hd__dfbbn_1_13/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_24 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_23/HI
+ sky130_fd_sc_hd__inv_1_32/Y FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__dfbbn_1_24/a_557_413# sky130_fd_sc_hd__dfbbn_1_24/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__dfbbn_1_24/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_581_47# sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# sky130_fd_sc_hd__dfbbn_1_24/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_35 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_37/HI
+ sky130_fd_sc_hd__inv_1_22/Y FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_35/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# sky130_fd_sc_hd__dfbbn_1_35/a_557_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_581_47# sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# sky130_fd_sc_hd__dfbbn_1_35/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_46 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_41/HI
+ sky130_fd_sc_hd__inv_1_50/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__dfbbn_1_46/a_557_413# sky130_fd_sc_hd__dfbbn_1_46/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_581_47# sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# sky130_fd_sc_hd__dfbbn_1_46/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_30 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_30/LO
+ sky130_fd_sc_hd__conb_1_30/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_41 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_41/LO
+ sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand3_1_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_20/Y
+ sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand3_1_0/a_193_47#
+ sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_29 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_18 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xtransmission_gate_3 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_123 V_GND sky130_fd_sc_hd__fill_4_194/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_101 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_112 V_GND sky130_fd_sc_hd__fill_4_215/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_134 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_145 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_156 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_167 V_GND sky130_fd_sc_hd__fill_4_320/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_29 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_29/Y sky130_fd_sc_hd__inv_16_29/A
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_18 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_16_19/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_14 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_16/HI
+ sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__dfbbn_1_14/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__dfbbn_1_14/a_557_413# sky130_fd_sc_hd__dfbbn_1_14/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_581_47# sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# sky130_fd_sc_hd__dfbbn_1_14/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_36 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_35/HI
+ sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__dfbbn_1_36/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__dfbbn_1_36/a_557_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# sky130_fd_sc_hd__dfbbn_1_36/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_47 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_39/HI
+ sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__dfbbn_1_47/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# sky130_fd_sc_hd__dfbbn_1_47/a_557_413# sky130_fd_sc_hd__dfbbn_1_47/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# sky130_fd_sc_hd__dfbbn_1_47/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_581_47# sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__dfbbn_1_47/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_25 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_24/HI
+ sky130_fd_sc_hd__inv_1_33/Y FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_25/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# sky130_fd_sc_hd__dfbbn_1_25/a_557_413# sky130_fd_sc_hd__dfbbn_1_25/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_581_47# sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# sky130_fd_sc_hd__dfbbn_1_25/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_31 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_31/LO
+ sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_20 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_20/LO
+ sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_42 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_42/LO
+ sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand3_1_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_66/Y
+ sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nand3_1_1/a_193_47#
+ sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_19 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xtransmission_gate_4 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_113 V_GND sky130_fd_sc_hd__fill_4_189/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_102 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_146 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_124 V_GND sky130_fd_sc_hd__fill_4_194/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_135 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_168 V_GND sky130_fd_sc_hd__fill_4_320/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_157 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_16_19 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_16_23/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__dfbbn_1_15 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_12/HI
+ sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# sky130_fd_sc_hd__dfbbn_1_15/a_557_413# sky130_fd_sc_hd__dfbbn_1_15/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__dfbbn_1_15/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_581_47# sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# sky130_fd_sc_hd__dfbbn_1_15/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_37 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_36/HI
+ sky130_fd_sc_hd__inv_1_43/Y RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_37/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# sky130_fd_sc_hd__dfbbn_1_37/a_557_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_581_47# sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# sky130_fd_sc_hd__dfbbn_1_37/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_48 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__dfbbn_1_48/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_43/HI
+ sky130_fd_sc_hd__inv_1_68/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_48/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# sky130_fd_sc_hd__dfbbn_1_48/a_557_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_381_47# sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_581_47# sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# sky130_fd_sc_hd__dfbbn_1_48/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_26 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_25/HI
+ sky130_fd_sc_hd__inv_1_30/Y FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__dfbbn_1_26/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# sky130_fd_sc_hd__dfbbn_1_26/a_557_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_581_47# sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# sky130_fd_sc_hd__dfbbn_1_26/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_10 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_10/LO
+ sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_21 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_21/LO
+ sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_32 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_32/LO
+ sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_43 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_43/LO
+ sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand3_1_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_51/Y
+ sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nand3_1_2/a_193_47#
+ sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__nand3_1
Xtransmission_gate_5 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_114 V_GND sky130_fd_sc_hd__fill_4_188/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_103 V_GND sky130_fd_sc_hd__fill_4_182/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_147 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_125 V_GND sky130_fd_sc_hd__fill_4_194/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_136 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_158 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_169 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_16 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_7/HI
+ sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_16/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# sky130_fd_sc_hd__dfbbn_1_16/a_557_413# sky130_fd_sc_hd__dfbbn_1_16/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_581_47# sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# sky130_fd_sc_hd__dfbbn_1_16/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_27 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_17/HI
+ sky130_fd_sc_hd__inv_1_26/Y RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__dfbbn_1_27/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__dfbbn_1_27/a_557_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_581_47# sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# sky130_fd_sc_hd__dfbbn_1_27/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_38 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_40/HI
+ sky130_fd_sc_hd__inv_1_55/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_38/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_38/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# sky130_fd_sc_hd__dfbbn_1_38/a_557_413# sky130_fd_sc_hd__dfbbn_1_38/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_38/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# sky130_fd_sc_hd__dfbbn_1_38/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_581_47# sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# sky130_fd_sc_hd__dfbbn_1_38/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__dfbbn_1_38/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_49 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_45/HI
+ sky130_fd_sc_hd__inv_1_61/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_49/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# sky130_fd_sc_hd__dfbbn_1_49/a_557_413# sky130_fd_sc_hd__dfbbn_1_49/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_581_47# sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# sky130_fd_sc_hd__dfbbn_1_49/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_11 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_11/LO
+ sky130_fd_sc_hd__conb_1_11/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_22 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_22/LO
+ sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_33 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_33/LO
+ sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_44 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_44/LO
+ sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1
Xtransmission_gate_6 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_104 V_GND sky130_fd_sc_hd__fill_4_184/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_115 V_GND sky130_fd_sc_hd__fill_4_189/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_126 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_137 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_159 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_148 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_28 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_32/HI
+ sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# sky130_fd_sc_hd__dfbbn_1_28/a_557_413# sky130_fd_sc_hd__dfbbn_1_28/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_581_47# sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# sky130_fd_sc_hd__dfbbn_1_28/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_17 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_19/HI
+ sky130_fd_sc_hd__inv_1_25/Y RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# sky130_fd_sc_hd__dfbbn_1_17/a_557_413# sky130_fd_sc_hd__dfbbn_1_17/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_581_47# sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# sky130_fd_sc_hd__dfbbn_1_17/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_39 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__dfbbn_1_39/Q_N sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_42/HI
+ sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_791_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# sky130_fd_sc_hd__dfbbn_1_39/a_557_413# sky130_fd_sc_hd__dfbbn_1_39/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_381_47# sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_581_47# sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# sky130_fd_sc_hd__dfbbn_1_39/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_12 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_12/LO
+ sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_34 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_34/LO
+ sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_45 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_45/LO
+ sky130_fd_sc_hd__conb_1_45/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_23 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_23/LO
+ sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1
Xtransmission_gate_7 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_105 V_GND sky130_fd_sc_hd__fill_4_182/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_116 V_GND sky130_fd_sc_hd__fill_4_188/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_138 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_127 V_GND sky130_fd_sc_hd__fill_4_215/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_149 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_18 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_21/HI
+ sky130_fd_sc_hd__inv_1_69/Y RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__dfbbn_1_18/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# sky130_fd_sc_hd__dfbbn_1_18/a_557_413# sky130_fd_sc_hd__dfbbn_1_18/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_581_47# sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# sky130_fd_sc_hd__dfbbn_1_18/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_29 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_31/HI
+ sky130_fd_sc_hd__inv_1_41/Y RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__dfbbn_1_29/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_791_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# sky130_fd_sc_hd__dfbbn_1_29/a_557_413# sky130_fd_sc_hd__dfbbn_1_29/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__dfbbn_1_29/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__dfbbn_1_29/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_581_47# sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# sky130_fd_sc_hd__dfbbn_1_29/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_13 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_13/LO
+ sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_35 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_35/LO
+ sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_24 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_24/LO
+ sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_46 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_46/LO
+ sky130_fd_sc_hd__conb_1_46/HI sky130_fd_sc_hd__conb_1
Xtransmission_gate_8 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_117 V_GND sky130_fd_sc_hd__fill_4_189/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_106 V_GND sky130_fd_sc_hd__fill_4_184/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_128 V_GND sky130_fd_sc_hd__fill_4_215/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_139 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_19 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_20/HI
+ sky130_fd_sc_hd__inv_1_28/Y RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__dfbbn_1_19/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# sky130_fd_sc_hd__dfbbn_1_19/a_557_413# sky130_fd_sc_hd__dfbbn_1_19/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_581_47# sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# sky130_fd_sc_hd__dfbbn_1_19/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_14 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_14/LO
+ sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_36 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_36/LO
+ sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_25 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_25/LO
+ sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_47 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_47/LO
+ sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__conb_1
Xtransmission_gate_9 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_118 V_GND sky130_fd_sc_hd__fill_4_188/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_129 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_107 V_GND sky130_fd_sc_hd__fill_4_215/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_15 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_15/LO
+ sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_37 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_37/LO
+ sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_26 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_26/LO
+ sky130_fd_sc_hd__conb_1_26/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_48 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_48/LO
+ sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_119 V_GND sky130_fd_sc_hd__fill_4_194/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_108 V_GND sky130_fd_sc_hd__fill_4_184/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_16 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_16/LO
+ sky130_fd_sc_hd__conb_1_16/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_38 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_38/LO
+ sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_27 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_27/LO
+ sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_49 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_49/LO
+ sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_109 V_GND sky130_fd_sc_hd__fill_4_182/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_28 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_28/LO
+ sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_17 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_17/LO
+ sky130_fd_sc_hd__conb_1_17/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_39 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_39/LO
+ sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_1/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_29 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_29/LO
+ sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_18 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_18/LO
+ sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_1_60 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__inv_1_60/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_2/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_19 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_19/LO
+ sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nand2_1_2/A
+ sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_50 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_61 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__conb_1_3/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_44/A
+ sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_40 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__inv_1_40/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_51 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_51/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_62 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__conb_1_4/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_8/A
+ sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_41 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_30 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__inv_1_30/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_52 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_52/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_63 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__inv_1_63/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_5/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__nand2_1_3/Y
+ sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfbbn_1_0 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_2/HI
+ sky130_fd_sc_hd__inv_1_4/Y FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_0/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_0/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# sky130_fd_sc_hd__dfbbn_1_0/a_557_413# sky130_fd_sc_hd__dfbbn_1_0/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_0/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__dfbbn_1_0/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_581_47# sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# sky130_fd_sc_hd__dfbbn_1_0/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# sky130_fd_sc_hd__dfbbn_1_0/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_42 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_42/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_20 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_20/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_31 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_64 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_64/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_53 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_53/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_6/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__nand2_8_9/A
+ sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__nand2_1
Xtransmission_gate_70 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__dfbbn_1_1 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_3/HI
+ sky130_fd_sc_hd__inv_1_2/Y FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__dfbbn_1_1/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__dfbbn_1_1/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# sky130_fd_sc_hd__dfbbn_1_1/a_557_413# sky130_fd_sc_hd__dfbbn_1_1/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_1/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# sky130_fd_sc_hd__dfbbn_1_1/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_581_47# sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# sky130_fd_sc_hd__dfbbn_1_1/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# sky130_fd_sc_hd__dfbbn_1_1/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_10 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_10/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_21 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_21/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_32 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_43 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_65 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_65/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_54 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_7/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__nand2_1_5/Y
+ sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__nand2_1
Xtransmission_gate_60 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_71 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__dfbbn_1_2 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_1/HI
+ sky130_fd_sc_hd__inv_1_0/Y FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_2/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_791_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_2/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# sky130_fd_sc_hd__dfbbn_1_2/a_557_413# sky130_fd_sc_hd__dfbbn_1_2/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__dfbbn_1_2/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# sky130_fd_sc_hd__dfbbn_1_2/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_581_47# sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# sky130_fd_sc_hd__dfbbn_1_2/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__dfbbn_1_2/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_0 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_0/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_11 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_11/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_22 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_22/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_33 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_44 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_2_0/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_66 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_66/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_55 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_0 V_GND V_HIGH V_GND V_HIGH transmission_gate_9/GN Reset
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_4_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__conb_1_8/HI
+ sky130_fd_sc_hd__conb_1
Xtransmission_gate_50 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_61 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_72 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__dfbbn_1_3 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_4/HI
+ sky130_fd_sc_hd__inv_1_1/Y FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_3/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_791_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__dfbbn_1_3/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_581_47# sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__dfbbn_1_3/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__dfbbn_1_3/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_1 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_1/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_12 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF16.Q
+ sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_23 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_23/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_45 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_34 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_67 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__inv_1_67/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_56 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_56/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_8/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_4_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__conb_1_9/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_8_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_19/Y sky130_fd_sc_hd__inv_1_23/A
+ sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_40 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_73 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_62 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_51 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__dfbbn_1_4 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_0/HI
+ sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_4/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# sky130_fd_sc_hd__dfbbn_1_4/a_557_413# sky130_fd_sc_hd__dfbbn_1_4/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__dfbbn_1_4/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# sky130_fd_sc_hd__dfbbn_1_4/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_581_47# sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# sky130_fd_sc_hd__dfbbn_1_4/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# sky130_fd_sc_hd__dfbbn_1_4/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_2 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_13 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF18.Q
+ sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_24 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_24/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_46 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_66/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_35 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__inv_1_35/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_57 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_68 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_16_4/Y
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_18/A
+ sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__nand2_8
Xtransmission_gate_41 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_30 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_52 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_74 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xtransmission_gate_63 Reset V_HIGH V_GND V_SENSE transmission_gate_9/GN transmission_gate
Xsky130_fd_sc_hd__dfbbn_1_5 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_9/HI
+ sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_5/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# sky130_fd_sc_hd__dfbbn_1_5/a_557_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_581_47# sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# sky130_fd_sc_hd__dfbbn_1_5/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# sky130_fd_sc_hd__dfbbn_1_5/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_3 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_3/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_14 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_36 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_47 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_47/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_25 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__inv_1_25/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_58 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__inv_1_58/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_69 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1
C0 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.352f
C1 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# V_LOW 0.0152f
C2 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.00182f
C3 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 5.79e-19
C4 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 7.35e-19
C5 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# -0.00282f
C6 V_SENSE sky130_fd_sc_hd__inv_1_68/Y 5.34e-19
C7 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_12/LO 1.65e-20
C8 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_19/A 0.00749f
C9 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_43/HI 5.38e-21
C10 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00134f
C11 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 8.05e-22
C12 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_16_41/Y 0.00278f
C13 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__nand3_1_2/Y 1.91e-19
C14 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__conb_1_4/HI -0.00677f
C15 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 7.37e-19
C16 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 5.16e-19
C17 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 9.96e-20
C18 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0.0116f
C19 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__conb_1_30/HI 8.47e-20
C20 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 3.13e-19
C21 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00382f
C22 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0.00128f
C23 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 5.09e-20
C24 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0199f
C25 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00374f
C26 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__conb_1_24/HI 4.02e-20
C27 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_381_47# -2.53e-20
C28 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 0.00108f
C29 sky130_fd_sc_hd__conb_1_42/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.223f
C30 sky130_fd_sc_hd__conb_1_2/LO RISING_COUNTER.COUNT_SUB_DFF1.Q 8.95e-21
C31 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_29/Y 0.0465f
C32 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_27_47# 0.0726f
C33 sky130_fd_sc_hd__conb_1_43/HI FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.438f
C34 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0.112f
C35 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# V_LOW 2.26e-20
C36 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__conb_1_10/HI 6.91e-19
C37 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# 7.02e-20
C38 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.2f
C39 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__conb_1_17/HI 0.023f
C40 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 0.00954f
C41 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 6.12e-19
C42 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 1.19e-19
C43 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00169f
C44 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_51/Y 0.506f
C45 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# sky130_fd_sc_hd__conb_1_38/HI 0.00183f
C46 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__conb_1_20/HI 0.0191f
C47 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__conb_1_46/HI 2.67e-20
C48 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_1_39/Y 4.43e-21
C49 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# V_LOW 3.56e-20
C50 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0251f
C51 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# -3.8e-20
C52 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# -0.00226f
C53 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.23e-20
C54 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# -1.76e-19
C55 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# -7.17e-20
C56 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_22/LO 0.00218f
C57 sky130_fd_sc_hd__conb_1_34/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 9.32e-21
C58 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.66e-21
C59 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# -0.0609f
C60 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 3.51e-21
C61 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_8/A 0.207f
C62 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 5.03e-20
C63 sky130_fd_sc_hd__dfbbn_1_33/a_581_47# sky130_fd_sc_hd__inv_1_34/Y 2.47e-19
C64 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 0.029f
C65 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_56/Y 9.73e-20
C66 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_6/HI 0.0116f
C67 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 3.23e-20
C68 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 2.02e-20
C69 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_26/Y -2.52e-19
C70 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# V_LOW -0.0127f
C71 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# 7.36e-19
C72 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# V_LOW 4.8e-20
C73 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_1_21/Y 0.00599f
C74 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0105f
C75 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_7/A 0.133f
C76 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_49/Y 2e-19
C77 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.22e-21
C78 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.44e-19
C79 sky130_fd_sc_hd__nand2_8_9/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 5.28e-20
C80 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__conb_1_51/HI 4.7e-20
C81 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 6.31e-19
C82 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__conb_1_12/HI -4.93e-19
C83 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# sky130_fd_sc_hd__conb_1_24/HI -6.57e-19
C84 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_44/A 0.00248f
C85 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00314f
C86 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__inv_1_38/Y 2.37e-21
C87 sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__inv_1_58/Y 0.00129f
C88 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 6.67e-19
C89 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 3.38e-20
C90 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 2.74e-20
C91 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# -1.61e-19
C92 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_473_413# -0.0122f
C93 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_46/A 0.00353f
C94 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__conb_1_10/HI 2.8e-19
C95 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# 4.57e-19
C96 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/Q_N -5.77e-19
C97 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 6.21e-20
C98 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 2.93e-20
C99 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__conb_1_29/HI 0.047f
C100 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00193f
C101 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_24/LO 6.71e-19
C102 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 0.00163f
C103 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__conb_1_2/HI 0.00138f
C104 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__inv_1_33/Y 7.14e-19
C105 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__inv_1_60/Y 4.33e-20
C106 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_44/HI 0.0272f
C107 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.00633f
C108 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__conb_1_43/HI 0.0234f
C109 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_45/Y 1.45e-19
C110 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_557_413# -3.67e-20
C111 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# -0.0242f
C112 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00294f
C113 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# Reset 0.00379f
C114 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# -0.00441f
C115 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__conb_1_28/HI 3.52e-20
C116 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 3.1e-21
C117 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# sky130_fd_sc_hd__conb_1_4/HI -9.33e-19
C118 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00201f
C119 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_24/Y 9.31e-19
C120 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 9.94e-19
C121 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 9.02e-20
C122 sky130_fd_sc_hd__inv_16_2/Y V_LOW 0.253f
C123 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 0.00175f
C124 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# -0.00117f
C125 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_381_47# -0.00832f
C126 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0222f
C127 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# -1.44e-20
C128 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 2.88e-21
C129 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.69e-21
C130 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00766f
C131 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_16_40/Y 0.0262f
C132 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00147f
C133 sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__conb_1_17/HI 0.00234f
C134 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.336f
C135 sky130_fd_sc_hd__conb_1_8/LO V_LOW 0.103f
C136 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -5.77e-20
C137 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# -2.52e-19
C138 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0.0581f
C139 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# V_LOW 0.0132f
C140 sky130_fd_sc_hd__inv_1_26/Y V_LOW 0.54f
C141 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# V_LOW 4.8e-20
C142 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 3.97e-20
C143 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__conb_1_46/HI 0.0045f
C144 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__conb_1_18/HI 6.57e-19
C145 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 2.12e-21
C146 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# V_LOW 0.00857f
C147 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_43/Y 7.51e-19
C148 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# -9.32e-20
C149 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__conb_1_5/HI 4.38e-20
C150 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_1_12/Y 0.00313f
C151 sky130_fd_sc_hd__inv_1_22/Y CLOCK_GEN.SR_Op.Q 6.45e-21
C152 sky130_fd_sc_hd__nand2_1_3/Y Reset 6.16e-19
C153 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.31e-19
C154 sky130_fd_sc_hd__inv_1_8/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 9.95e-19
C155 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.06e-20
C156 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 1.2e-19
C157 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# V_LOW 0.0459f
C158 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0529f
C159 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 2.01e-19
C160 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__inv_1_26/Y 0.00222f
C161 sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# V_LOW -6.55e-19
C162 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0.01f
C163 sky130_fd_sc_hd__inv_1_52/A CLOCK_GEN.SR_Op.Q 0.00325f
C164 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__inv_1_7/Y 4.76e-20
C165 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 6.04e-20
C166 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 9.24e-20
C167 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 3.29e-21
C168 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_24/HI 1.48e-22
C169 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 3.09e-19
C170 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_24/A 1.22e-19
C171 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__conb_1_12/HI -1.15e-19
C172 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.69e-19
C173 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0455f
C174 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__inv_1_12/Y 2.51e-20
C175 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__conb_1_32/HI 9.8e-19
C176 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 0.00359f
C177 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# V_LOW 0.013f
C178 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# -2.57e-20
C179 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_12/Y 0.141f
C180 sky130_fd_sc_hd__inv_16_51/Y CLOCK_GEN.SR_Op.Q 0.0194f
C181 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 9.75e-19
C182 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 1.68e-19
C183 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 2.52e-19
C184 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__conb_1_10/HI 2.43e-19
C185 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00143f
C186 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_29/HI 0.00668f
C187 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 0.0012f
C188 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.28e-21
C189 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_19/Y 0.121f
C190 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__conb_1_26/HI 0.00369f
C191 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0.0266f
C192 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 9.67e-22
C193 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__conb_1_28/HI 7.28e-20
C194 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_49/A 0.29f
C195 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__inv_1_50/Y 0.0102f
C196 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__conb_1_4/HI 0.00347f
C197 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 1.05e-19
C198 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 8.23e-19
C199 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 1.11e-20
C200 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# -0.00133f
C201 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# -0.00832f
C202 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# sky130_fd_sc_hd__conb_1_44/HI 2.22e-20
C203 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# 4.31e-19
C204 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0247f
C205 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# Reset 2.71e-19
C206 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# -0.00148f
C207 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 3.16e-21
C208 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_16_40/Y 2.33e-21
C209 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# CLOCK_GEN.SR_Op.Q 5.75e-20
C210 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__conb_1_4/HI 4.11e-19
C211 sky130_fd_sc_hd__dfbbn_1_51/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0121f
C212 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00287f
C213 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# sky130_fd_sc_hd__inv_16_42/Y 0.00106f
C214 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/Q_N 2.78e-19
C215 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 5.77e-19
C216 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0296f
C217 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 2.43e-20
C218 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_381_47# 0.00105f
C219 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.169f
C220 sky130_fd_sc_hd__fill_4_189/VPB V_LOW 0.854f
C221 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00124f
C222 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__inv_1_35/Y 1.79e-19
C223 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0.03f
C224 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 3.21e-21
C225 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0399f
C226 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.204f
C227 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_557_413# -3.67e-20
C228 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# -0.00623f
C229 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.36e-19
C230 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00105f
C231 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# -1.76e-19
C232 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# 3.94e-21
C233 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_473_413# -3.86e-20
C234 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_941_21# -1.61e-20
C235 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# sky130_fd_sc_hd__conb_1_46/HI -0.00262f
C236 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# sky130_fd_sc_hd__conb_1_18/HI -2.65e-20
C237 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0024f
C238 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__conb_1_24/HI 0.0122f
C239 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 4.4e-19
C240 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.327f
C241 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_1_40/Y 3.7e-19
C242 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/Q_N -4.78e-20
C243 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# sky130_fd_sc_hd__conb_1_5/HI 7.59e-20
C244 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__conb_1_9/LO 0.0401f
C245 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_22/Y 7.36e-20
C246 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_32/Y 0.0219f
C247 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -1.67e-19
C248 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -9.88e-20
C249 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_381_47# -4.37e-20
C250 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__inv_1_29/Y 1.98e-19
C251 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 4.5e-20
C252 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.67e-20
C253 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# V_LOW 2.94e-20
C254 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00147f
C255 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__inv_1_49/Y 2.48e-19
C256 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_32/HI 5.37e-20
C257 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_5/HI -0.00181f
C258 sky130_fd_sc_hd__inv_1_46/A CLOCK_GEN.SR_Op.Q 0.162f
C259 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_7/HI 2.2e-19
C260 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__inv_1_40/Y 2.64e-20
C261 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.35e-19
C262 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__conb_1_10/LO 1.3e-20
C263 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.21e-19
C264 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.27e-20
C265 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_66/Y 3.02e-20
C266 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__conb_1_19/HI 8.1e-20
C267 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00161f
C268 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_48/A 0.00994f
C269 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_1_44/A 0.00366f
C270 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00312f
C271 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.55e-19
C272 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__inv_1_12/Y 1.06e-19
C273 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_26/Y 0.382f
C274 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__inv_1_13/Y 6.12e-20
C275 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.45e-21
C276 sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# sky130_fd_sc_hd__conb_1_32/HI 0.00196f
C277 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 0.00433f
C278 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 8.84e-20
C279 sky130_fd_sc_hd__conb_1_9/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 1.38e-21
C280 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 4.71e-20
C281 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 2.01e-20
C282 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# -4.66e-20
C283 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__conb_1_25/HI 7.4e-20
C284 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/Q_N 7.56e-19
C285 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 6.4e-20
C286 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# 1.44e-19
C287 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_1_13/Y 0.0139f
C288 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 8.17e-19
C289 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_67/A 0.00392f
C290 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_791_47# 0.00616f
C291 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_35/Y 0.201f
C292 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_33/Y 4.43e-21
C293 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__conb_1_21/HI 0.00191f
C294 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# V_LOW 0.0114f
C295 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 1.31e-20
C296 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 1.81e-19
C297 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_10/Y 3.71e-19
C298 RISING_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 8.03e-21
C299 FULL_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0238f
C300 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# V_LOW 3.56e-20
C301 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0211f
C302 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 0.0298f
C303 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_56/A 6.08e-21
C304 sky130_fd_sc_hd__inv_1_0/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 2.95e-19
C305 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00386f
C306 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_19/A 0.00226f
C307 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_3/Y 1.93e-20
C308 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# V_LOW -0.00389f
C309 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_48/A 3.03e-19
C310 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_1_27/Y 0.00166f
C311 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 0.0116f
C312 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.81e-20
C313 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 7.04e-19
C314 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0717f
C315 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.07e-20
C316 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 1.54e-19
C317 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.67e-20
C318 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 6.04e-19
C319 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_44/A 7.75e-22
C320 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# -6.57e-19
C321 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 1.54e-19
C322 FULL_COUNTER.COUNT_SUB_DFF14.Q V_LOW 1.92f
C323 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00276f
C324 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# V_LOW 0.0338f
C325 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__conb_1_33/HI -0.00889f
C326 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/Q_N 4.55e-20
C327 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nor2_1_0/Y 0.00422f
C328 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.0461f
C329 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00304f
C330 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_37/Q_N 1.29e-19
C331 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_647_21# 1.74e-20
C332 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 0.00194f
C333 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_891_329# -0.00159f
C334 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# -0.0085f
C335 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.75e-20
C336 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 9.88e-22
C337 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__inv_1_69/Y 0.00318f
C338 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_19/A 0.0434f
C339 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# -2.57e-20
C340 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.86e-21
C341 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_4/Y 0.0036f
C342 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.149f
C343 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_11/HI 0.00248f
C344 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_58/Y 1.71e-19
C345 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.34e-19
C346 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# V_LOW 0.00545f
C347 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 7e-19
C348 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_42/Y 0.198f
C349 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__inv_1_40/Y 7.6e-19
C350 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.167f
C351 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__conb_1_26/HI 5.87e-20
C352 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 0.00483f
C353 sky130_fd_sc_hd__inv_1_54/Y V_LOW 0.217f
C354 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__conb_1_21/HI 2.57e-21
C355 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__conb_1_28/HI 5.83e-19
C356 sky130_fd_sc_hd__inv_1_16/Y V_LOW 0.403f
C357 sky130_fd_sc_hd__inv_1_24/A CLOCK_GEN.SR_Op.Q 0.0266f
C358 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.36e-19
C359 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__nand2_1_3/Y 3.02e-21
C360 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__inv_1_25/Y 7.18e-21
C361 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_473_413# 0.0344f
C362 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_19/LO 0.00178f
C363 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# sky130_fd_sc_hd__conb_1_32/HI 8.74e-19
C364 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_1_61/Y 1.22e-19
C365 sky130_fd_sc_hd__conb_1_0/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0283f
C366 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.28e-20
C367 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00882f
C368 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__inv_1_38/Y 6.24e-19
C369 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_20/HI 7.29e-19
C370 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_45/A 0.0767f
C371 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 2.78e-21
C372 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__nand2_8_8/A 0.00288f
C373 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.02e-21
C374 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__conb_1_19/HI 2.73e-20
C375 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__inv_1_44/A 4.7e-19
C376 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__conb_1_23/HI 0.0017f
C377 sky130_fd_sc_hd__dfbbn_1_39/Q_N FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0253f
C378 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 3.19e-20
C379 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.5e-19
C380 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# -0.0158f
C381 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# -9.34e-19
C382 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_791_47# 4.97e-19
C383 sky130_fd_sc_hd__inv_16_41/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.14f
C384 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__conb_1_3/HI 0.00262f
C385 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# -0.00115f
C386 V_SENSE sky130_fd_sc_hd__inv_16_49/Y 2.48f
C387 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__nand2_1_2/A 0.00147f
C388 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_30/HI 0.0354f
C389 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__conb_1_46/LO 0.0117f
C390 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 2.19e-19
C391 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__conb_1_25/HI 1.69e-19
C392 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0513f
C393 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 7.41e-19
C394 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# 4.18e-19
C395 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__inv_1_13/Y 0.0432f
C396 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_1_39/Y 1.32e-21
C397 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.13e-19
C398 sky130_fd_sc_hd__inv_1_41/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.466f
C399 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_1_31/Y 9.34e-19
C400 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__conb_1_21/HI 1.35e-20
C401 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/Q_N -9.56e-20
C402 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI -2.03e-20
C403 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_16/LO 0.0148f
C404 sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__inv_1_53/Y 1.82e-19
C405 sky130_fd_sc_hd__conb_1_34/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 5.88e-20
C406 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 4.38e-19
C407 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0283f
C408 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__inv_1_45/Y 0.00222f
C409 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.22e-21
C410 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__conb_1_11/HI 0.00317f
C411 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 0.00366f
C412 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 4.2e-19
C413 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 8.46e-19
C414 sky130_fd_sc_hd__conb_1_8/HI V_LOW 0.152f
C415 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0205f
C416 sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00161f
C417 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0117f
C418 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0422f
C419 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__inv_1_10/Y 0.0374f
C420 sky130_fd_sc_hd__nand2_8_9/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 7.84e-21
C421 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_48/Y 1.61e-20
C422 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_56/Y 1.15e-19
C423 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# V_LOW 4.8e-20
C424 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# -5.54e-21
C425 sky130_fd_sc_hd__inv_1_2/Y V_LOW 0.207f
C426 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# V_LOW 0.0151f
C427 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_557_413# 7.19e-19
C428 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# sky130_fd_sc_hd__conb_1_33/HI -9.57e-19
C429 sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.00525f
C430 sky130_fd_sc_hd__inv_1_57/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00579f
C431 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__nand2_8_4/Y 0.00158f
C432 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__conb_1_7/HI 7.71e-21
C433 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# -0.00196f
C434 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_4/LO 0.00305f
C435 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# sky130_fd_sc_hd__conb_1_31/HI -6.57e-19
C436 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# sky130_fd_sc_hd__inv_1_69/Y 1.07e-21
C437 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__inv_1_13/Y 2.45e-19
C438 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__conb_1_11/LO 9.17e-19
C439 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_1_41/Y 1.26e-19
C440 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 8.11e-19
C441 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.89e-19
C442 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# V_LOW -2.78e-35
C443 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 9.76e-20
C444 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# -4.66e-20
C445 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_381_47# -3.79e-20
C446 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 5.43e-19
C447 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 7.46e-20
C448 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/Q_N -9.56e-20
C449 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.86e-21
C450 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00878f
C451 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00227f
C452 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# 0.00501f
C453 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.18e-19
C454 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_19/Y 3.38e-19
C455 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 4.54e-20
C456 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_66/A 0.106f
C457 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_47/Y 0.00212f
C458 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__conb_1_2/HI 0.0303f
C459 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# V_LOW 0.0416f
C460 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 2.81e-19
C461 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 3.61e-19
C462 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 9.26e-19
C463 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.235f
C464 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# V_LOW 0.00458f
C465 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# Reset 0.00457f
C466 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.17f
C467 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_51/Y 0.00145f
C468 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__conb_1_23/HI -0.0127f
C469 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__conb_1_45/LO 2.32e-20
C470 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 1.58e-19
C471 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__inv_1_1/Y 0.00466f
C472 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# -6.8e-19
C473 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.33e-19
C474 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# 9.42e-20
C475 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# sky130_fd_sc_hd__conb_1_3/HI 1.15e-21
C476 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00332f
C477 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_581_47# -7.91e-19
C478 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_59/Y 0.194f
C479 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_1_60/Y 3.31e-20
C480 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# sky130_fd_sc_hd__conb_1_30/HI 9.52e-19
C481 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# -1.24e-20
C482 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__conb_1_25/HI 0.00116f
C483 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.056f
C484 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 5.13e-19
C485 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# V_LOW 0.0177f
C486 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__inv_1_14/Y 1.72e-20
C487 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_17/a_557_413# 3.74e-20
C488 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.105f
C489 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__conb_1_45/HI -2.07e-19
C490 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__conb_1_41/HI 0.00478f
C491 sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF12.Q 0.128f
C492 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand3_1_2/Y 4.49e-21
C493 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_66/A 5.43e-20
C494 sky130_fd_sc_hd__inv_1_42/Y Reset 0.00435f
C495 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_6/LO 1.69e-20
C496 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.92e-21
C497 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.19e-19
C498 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# sky130_fd_sc_hd__conb_1_11/HI 1.15e-20
C499 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_66/A 0.0755f
C500 sky130_fd_sc_hd__dfbbn_1_13/Q_N FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0166f
C501 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_10/LO 3.51e-20
C502 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_38/HI 1.15e-20
C503 V_SENSE RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0671f
C504 sky130_fd_sc_hd__conb_1_6/LO V_LOW 0.0879f
C505 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.81e-19
C506 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# -0.054f
C507 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# 3.58e-20
C508 sky130_fd_sc_hd__inv_16_2/Y V_HIGH 0.693f
C509 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 7.48e-19
C510 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 9.68e-20
C511 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 1.2e-19
C512 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_47/HI 0.0851f
C513 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__conb_1_33/HI -2.17e-19
C514 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_19/A 0.00764f
C515 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 0.00999f
C516 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__inv_1_28/Y 0.0103f
C517 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__inv_2_0/A 0.00623f
C518 sky130_fd_sc_hd__inv_16_20/A sky130_fd_sc_hd__inv_16_24/Y 0.0442f
C519 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_1_21/Y 0.0157f
C520 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# -0.00263f
C521 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# -5.54e-21
C522 sky130_fd_sc_hd__conb_1_5/LO FULL_COUNTER.COUNT_SUB_DFF6.Q 4.41e-20
C523 sky130_fd_sc_hd__dfbbn_1_50/Q_N V_LOW -2.68e-19
C524 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 1.5e-19
C525 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_41/Y 0.645f
C526 sky130_fd_sc_hd__inv_16_15/Y sky130_fd_sc_hd__inv_16_8/A 9.54e-22
C527 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_56/Y 0.0742f
C528 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_473_413# -0.012f
C529 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -0.00966f
C530 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.31e-20
C531 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 2.83e-20
C532 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 5.52e-21
C533 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__inv_1_55/Y 0.0292f
C534 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_67/A 2.05e-21
C535 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__conb_1_2/HI 0.0517f
C536 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# V_LOW 2.94e-20
C537 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 0.0021f
C538 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# 7.25e-19
C539 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.47e-21
C540 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# V_LOW -0.323f
C541 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 5.08e-20
C542 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_39/HI 2.05e-19
C543 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# CLOCK_GEN.SR_Op.Q 8.98e-19
C544 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# -8.61e-20
C545 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# V_LOW 4.8e-20
C546 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_16_19/Y 3.23e-19
C547 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0242f
C548 sky130_fd_sc_hd__conb_1_3/LO V_LOW 0.0429f
C549 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 2.82e-19
C550 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_6/Y 0.0728f
C551 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00501f
C552 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# V_LOW -0.311f
C553 sky130_fd_sc_hd__dfbbn_1_37/Q_N FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00404f
C554 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 1.43e-19
C555 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00129f
C556 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00626f
C557 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 7.28e-20
C558 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0398f
C559 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__conb_1_9/HI 4.46e-19
C560 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 2.33e-20
C561 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_581_47# -2.6e-20
C562 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 8.84e-20
C563 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.114f
C564 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_1_39/Y 3.79e-20
C565 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# V_LOW 0.00105f
C566 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__inv_1_39/Y 8.76e-19
C567 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 0.00174f
C568 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_1_8/Y 2.55e-21
C569 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__nand3_1_1/Y 0.00891f
C570 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_1_44/A 0.0518f
C571 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# sky130_fd_sc_hd__conb_1_41/HI -0.00262f
C572 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 0.00773f
C573 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_23/A 4.49e-19
C574 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_47/Y 2.14e-21
C575 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 7.91e-19
C576 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__conb_1_4/HI 5.89e-19
C577 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 4.59e-21
C578 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__inv_1_38/Y 0.00491f
C579 V_SENSE sky130_fd_sc_hd__conb_1_43/HI 4.83e-19
C580 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00143f
C581 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__conb_1_16/LO 5.37e-20
C582 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0188f
C583 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_1_32/Y 1.07e-19
C584 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00337f
C585 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/Q_N -4.33e-20
C586 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_65/A 9.19e-20
C587 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__conb_1_47/HI 2.04e-19
C588 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0385f
C589 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 6.31e-21
C590 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 3.23e-21
C591 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__conb_1_51/HI -3.44e-19
C592 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.76e-19
C593 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 0.245f
C594 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# -0.00834f
C595 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -1.61e-19
C596 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 1.95e-19
C597 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 1.79e-19
C598 sky130_fd_sc_hd__conb_1_0/LO V_LOW 0.0909f
C599 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# sky130_fd_sc_hd__inv_1_44/A 1.99e-19
C600 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_8_8/A 3.04e-20
C601 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# -9.32e-20
C602 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# V_LOW 0.0422f
C603 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0223f
C604 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_31/Q_N -3.55e-33
C605 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__conb_1_6/HI 0.00731f
C606 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 2.31e-19
C607 FULL_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0194f
C608 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.0407f
C609 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# -2.57e-20
C610 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0023f
C611 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00865f
C612 sky130_fd_sc_hd__inv_1_0/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 2.15e-20
C613 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_58/Y 0.00263f
C614 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__inv_1_47/A 0.00311f
C615 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__inv_1_28/Y 0.244f
C616 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__conb_1_15/HI 0.00135f
C617 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_55/Y 0.357f
C618 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 0.00147f
C619 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__conb_1_8/HI -0.00218f
C620 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -2.6e-19
C621 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# -3.48e-19
C622 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 8e-21
C623 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 3.67e-21
C624 sky130_fd_sc_hd__dfbbn_1_15/Q_N V_LOW -0.00504f
C625 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# V_LOW -0.0819f
C626 FULL_COUNTER.COUNT_SUB_DFF13.Q V_LOW 2.03f
C627 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_44/A 0.01f
C628 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_581_47# -7.91e-19
C629 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__inv_1_13/Y 0.1f
C630 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# V_LOW -0.00446f
C631 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00161f
C632 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# V_LOW 2.26e-20
C633 V_SENSE sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 1.15e-19
C634 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__conb_1_45/LO 1.2e-19
C635 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0278f
C636 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF18.Q 0.427f
C637 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_10/Y 8.35e-20
C638 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF0.Q 8.28e-19
C639 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_7/HI -0.00266f
C640 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# V_LOW 0.0153f
C641 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__conb_1_20/HI 1.55e-19
C642 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.0327f
C643 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# V_LOW -9.15e-19
C644 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_7/HI 0.0768f
C645 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.74e-19
C646 V_SENSE FULL_COUNTER.COUNT_SUB_DFF1.Q 0.117f
C647 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# 5.49e-19
C648 sky130_fd_sc_hd__dfbbn_1_32/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 7.04e-20
C649 CLOCK_GEN.SR_Op.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00175f
C650 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__dfbbn_1_0/a_193_47# 2.19e-19
C651 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_42/Y 3.19e-19
C652 sky130_fd_sc_hd__conb_1_0/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0258f
C653 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 0.00221f
C654 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# V_LOW -3.04e-19
C655 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# V_LOW 2.26e-20
C656 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/Q_N 4.8e-19
C657 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.78e-21
C658 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_8/A 2.88e-19
C659 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 7.35e-19
C660 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.09e-19
C661 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.55e-20
C662 sky130_fd_sc_hd__conb_1_12/HI FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0301f
C663 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_67/A 0.439f
C664 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_16_24/Y 7.43e-20
C665 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0198f
C666 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0313f
C667 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_40/Y 6e-19
C668 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# -2.57e-20
C669 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0502f
C670 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/Q_N -4.78e-20
C671 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 0.0398f
C672 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# V_LOW -6.55e-19
C673 sky130_fd_sc_hd__inv_16_49/Y CLOCK_GEN.SR_Op.Q 0.0207f
C674 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 0.0353f
C675 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 3.75e-19
C676 sky130_fd_sc_hd__conb_1_16/HI V_LOW 0.0139f
C677 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 6.72e-20
C678 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 6.72e-20
C679 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.21e-19
C680 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 1.37e-20
C681 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 2.76e-20
C682 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0209f
C683 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# sky130_fd_sc_hd__conb_1_15/HI -2.65e-20
C684 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF15.Q 4.76e-19
C685 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 9.03e-20
C686 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 0.00484f
C687 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# sky130_fd_sc_hd__conb_1_8/HI -0.00116f
C688 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 8.17e-19
C689 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_2_0/A 9.7e-21
C690 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -6.22e-19
C691 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# -0.00449f
C692 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# -6.23e-21
C693 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 6.4e-21
C694 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# V_LOW -2.68e-19
C695 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_381_47# 0.00286f
C696 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/Q_N 7.72e-21
C697 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_28/HI 2.23e-20
C698 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_48/Y 9.73e-19
C699 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 0.00109f
C700 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# -2.52e-19
C701 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# -0.00144f
C702 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__conb_1_7/HI -2.07e-19
C703 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00211f
C704 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 0.00841f
C705 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.556f
C706 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__conb_1_0/HI 5.75e-20
C707 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__nand3_1_1/Y 0.00384f
C708 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00288f
C709 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 0.027f
C710 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.37e-21
C711 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.65e-21
C712 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# sky130_fd_sc_hd__inv_1_13/Y 1.14e-20
C713 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_50/HI -8.38e-19
C714 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# -0.00125f
C715 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -6.22e-19
C716 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# -4.37e-20
C717 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0227f
C718 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# -0.187f
C719 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_581_47# 6.42e-19
C720 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_53/A 1.38e-20
C721 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_1_22/Y 4.5e-20
C722 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_38/HI 0.00307f
C723 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.62e-21
C724 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 3.23e-19
C725 sky130_fd_sc_hd__inv_1_35/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 7.73e-20
C726 sky130_fd_sc_hd__inv_1_58/Y sky130_fd_sc_hd__inv_1_30/Y 0.0406f
C727 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# V_LOW -0.00266f
C728 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_25/HI 0.358f
C729 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.55e-19
C730 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 7.18e-19
C731 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand3_1_2/a_109_47# 2.15e-19
C732 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.00267f
C733 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00482f
C734 sky130_fd_sc_hd__inv_1_3/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0219f
C735 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0571f
C736 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_25/Y 5.18e-20
C737 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 9.85e-19
C738 sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.199f
C739 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 6.87e-20
C740 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 1.45e-19
C741 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 6.87e-20
C742 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 0.0126f
C743 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 1.45e-19
C744 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0.0128f
C745 sky130_fd_sc_hd__inv_1_28/Y V_LOW 0.191f
C746 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 0.00446f
C747 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_473_413# -0.00312f
C748 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_647_21# -0.00122f
C749 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.68e-19
C750 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_0/Y 0.0574f
C751 FALLING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 8.17e-19
C752 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# V_LOW -0.00389f
C753 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.11f
C754 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 2e-19
C755 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# -5.54e-21
C756 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# -0.00138f
C757 sky130_fd_sc_hd__conb_1_46/HI FALLING_COUNTER.COUNT_SUB_DFF6.Q 5.13e-20
C758 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_16_2/Y 0.153f
C759 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__nor2_1_0/Y 1.21e-19
C760 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_791_47# 9.79e-21
C761 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/Q_N -4.78e-20
C762 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 1.88e-20
C763 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 1.69e-20
C764 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__conb_1_35/HI -0.0026f
C765 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_66/Y 1.13e-20
C766 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 2.72e-21
C767 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.3e-20
C768 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__conb_1_40/HI 0.004f
C769 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 1.79e-19
C770 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_647_21# 1.97e-20
C771 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__conb_1_46/HI 5.42e-19
C772 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00222f
C773 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# V_LOW -0.00751f
C774 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# V_LOW 3.56e-20
C775 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 0.00942f
C776 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_381_47# -2.53e-20
C777 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# -5.16e-20
C778 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# -1.76e-19
C779 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 1.68e-19
C780 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 2.52e-19
C781 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 9.75e-19
C782 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.088f
C783 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_48/Y 0.00387f
C784 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_37/HI 0.86f
C785 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00111f
C786 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_39/HI 9.87e-21
C787 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 9.52e-20
C788 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 9.52e-20
C789 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 0.00152f
C790 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 5.17e-20
C791 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 5.37e-19
C792 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 2.96e-19
C793 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_56/A 0.00152f
C794 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__inv_1_26/Y 7.64e-20
C795 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# FULL_COUNTER.COUNT_SUB_DFF12.Q 9.76e-19
C796 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0233f
C797 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_47/Y 0.00817f
C798 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 6.05e-21
C799 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 7.72e-20
C800 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.88e-20
C801 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.138f
C802 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__conb_1_27/HI 0.00329f
C803 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.72e-20
C804 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.93e-19
C805 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# V_LOW 0.00117f
C806 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__conb_1_50/HI -0.00575f
C807 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__conb_1_9/HI 4.47e-20
C808 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0311f
C809 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_46/A 0.236f
C810 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.48e-21
C811 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00343f
C812 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.04e-20
C813 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_13/LO 1.33e-19
C814 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0253f
C815 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_4/LO 4.26e-19
C816 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_47/Y 3.77e-22
C817 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.94e-21
C818 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.0701f
C819 sky130_fd_sc_hd__dfbbn_1_44/a_581_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 7.59e-20
C820 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__conb_1_14/HI 0.00488f
C821 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0355f
C822 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__conb_1_11/HI 4.58e-20
C823 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 0.00118f
C824 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 4.87e-21
C825 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 7.77e-19
C826 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 8.54e-21
C827 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.08e-20
C828 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__conb_1_29/HI 0.0414f
C829 sky130_fd_sc_hd__inv_1_15/Y V_LOW 0.441f
C830 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_39/HI -0.00195f
C831 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_27/Y 0.00332f
C832 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.00379f
C833 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_56/A 0.00574f
C834 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 0.00275f
C835 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__inv_1_50/Y 7.22e-21
C836 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_33/HI 4.84e-21
C837 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0323f
C838 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 5.66e-19
C839 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/Q_N 5.66e-19
C840 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_31/HI 0.0183f
C841 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_33/Y 4.36e-19
C842 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.9e-20
C843 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__inv_1_0/Y 3.94e-21
C844 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0193f
C845 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 6.69e-19
C846 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# -9.32e-20
C847 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_19/Y 0.0201f
C848 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__inv_1_59/Y 0.0446f
C849 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 8.02e-21
C850 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 2.66e-21
C851 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.19e-19
C852 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.92e-20
C853 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.0313f
C854 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# V_LOW 2.94e-20
C855 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# -0.00631f
C856 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# -0.00988f
C857 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -0.00126f
C858 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# -2.37e-19
C859 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__inv_1_49/Y 2.47e-20
C860 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 0.00837f
C861 V_SENSE sky130_fd_sc_hd__inv_16_55/Y 0.358f
C862 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 2.06e-20
C863 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00306f
C864 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# -0.00141f
C865 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 1.62e-20
C866 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_40/LO 7.93e-20
C867 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 2.01e-20
C868 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 4.71e-20
C869 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 0.0395f
C870 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_193_47# -0.2f
C871 sky130_fd_sc_hd__conb_1_1/HI V_LOW 0.159f
C872 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.023f
C873 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0021f
C874 sky130_fd_sc_hd__inv_1_6/Y V_LOW 0.144f
C875 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 0.0021f
C876 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 2.07e-19
C877 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 0.0114f
C878 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_791_47# 1.68e-19
C879 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 3.12e-20
C880 FULL_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0314f
C881 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0518f
C882 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 8.74e-20
C883 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# sky130_fd_sc_hd__inv_1_2/Y 7.97e-21
C884 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 4.54e-21
C885 sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__conb_1_19/HI 0.00607f
C886 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# V_LOW 3.56e-20
C887 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_24/A 0.0019f
C888 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# 8.69e-19
C889 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_29/HI 1.64e-19
C890 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 0.00198f
C891 sky130_fd_sc_hd__inv_1_68/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.42e-20
C892 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# -3.79e-20
C893 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# -4.66e-20
C894 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.2e-19
C895 sky130_fd_sc_hd__inv_16_6/A FULL_COUNTER.COUNT_SUB_DFF2.Q 0.325f
C896 sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# sky130_fd_sc_hd__conb_1_9/HI -2.65e-20
C897 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/Q_N -9.56e-20
C898 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__conb_1_4/HI 0.00456f
C899 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00259f
C900 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# V_LOW 0.00694f
C901 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.0593f
C902 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 4.21e-19
C903 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0128f
C904 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# sky130_fd_sc_hd__conb_1_14/HI 1.68e-19
C905 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 4.2e-19
C906 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_67/A 0.519f
C907 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_21/Y 0.139f
C908 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0214f
C909 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.04f
C910 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 4.55e-19
C911 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 8.96e-19
C912 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 1.86e-20
C913 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 1.12e-20
C914 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_38/Y 9.87e-21
C915 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__conb_1_39/HI -2.07e-19
C916 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_381_47# 9.87e-20
C917 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 3.46e-20
C918 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00463f
C919 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# sky130_fd_sc_hd__inv_1_50/Y 2.78e-22
C920 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00287f
C921 V_SENSE FULL_COUNTER.COUNT_SUB_DFF0.Q 0.169f
C922 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.223f
C923 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 7.79e-21
C924 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_8/LO 0.00128f
C925 sky130_fd_sc_hd__conb_1_41/HI V_LOW 0.177f
C926 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_27/Y 0.0712f
C927 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# Reset 8.68e-19
C928 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_891_329# 6.63e-21
C929 CLOCK_GEN.SR_Op.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 4.05e-19
C930 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_1/Y 0.0372f
C931 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 1.96e-20
C932 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 6.14e-20
C933 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 2.3e-21
C934 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.53e-20
C935 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0807f
C936 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 8.97e-19
C937 sky130_fd_sc_hd__conb_1_0/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.956f
C938 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/Q_N -4.33e-20
C939 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# sky130_fd_sc_hd__conb_1_2/HI 5.79e-19
C940 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_66/A 1.12e-19
C941 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00954f
C942 sky130_fd_sc_hd__conb_1_27/LO RISING_COUNTER.COUNT_SUB_DFF4.Q 1.31e-20
C943 sky130_fd_sc_hd__inv_1_65/A V_LOW 0.412f
C944 sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_32/Y 0.0115f
C945 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# -0.00519f
C946 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_26/Y 3.78e-20
C947 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.01e-19
C948 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# -0.2f
C949 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.53e-20
C950 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_25/HI 9.64e-21
C951 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.38e-19
C952 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_12/LO 1.82e-19
C953 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 0.0074f
C954 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_15/HI 4.84e-20
C955 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 2.97e-19
C956 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__inv_1_1/Y 1.12e-20
C957 sky130_fd_sc_hd__conb_1_36/HI V_LOW 0.197f
C958 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# -1.66e-19
C959 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 1.47e-21
C960 sky130_fd_sc_hd__inv_1_67/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 1.41e-19
C961 sky130_fd_sc_hd__inv_1_25/Y sky130_fd_sc_hd__inv_1_26/Y 0.0227f
C962 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__inv_1_40/Y 9.13e-21
C963 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_1_19/A 1.67e-19
C964 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 7.89e-21
C965 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_16_19/Y 1.38e-20
C966 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.42e-19
C967 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.13e-19
C968 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_40/a_941_21# 1.68e-19
C969 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0039f
C970 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 7.97e-20
C971 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__conb_1_17/HI 0.00364f
C972 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 5.1e-20
C973 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_791_47# 6.99e-20
C974 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 2.01e-20
C975 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0249f
C976 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0119f
C977 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.29e-22
C978 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 2.07e-19
C979 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 8.34e-19
C980 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 8.22e-19
C981 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.18e-21
C982 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.57e-20
C983 V_SENSE sky130_fd_sc_hd__inv_16_44/Y 1.96f
C984 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0199f
C985 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 1.74e-20
C986 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 0.00181f
C987 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 6.87e-22
C988 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# -3.06e-20
C989 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# -6.43e-20
C990 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__conb_1_39/HI 0.0225f
C991 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__inv_1_66/A 5.04e-19
C992 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 1.8e-20
C993 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# V_LOW -8.72e-19
C994 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# V_LOW -0.313f
C995 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# V_LOW 2.26e-20
C996 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_891_329# -2.2e-20
C997 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# -4.1e-19
C998 sky130_fd_sc_hd__dfbbn_1_19/Q_N V_LOW -0.00253f
C999 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.41e-21
C1000 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# V_LOW 0.042f
C1001 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__nand2_8_1/a_27_47# 0.0032f
C1002 sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# sky130_fd_sc_hd__conb_1_3/HI -6.57e-19
C1003 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# sky130_fd_sc_hd__inv_1_60/Y 8.64e-19
C1004 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.0306f
C1005 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0156f
C1006 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_16_2/Y 9.59e-20
C1007 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# -4.66e-20
C1008 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 0.00153f
C1009 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00224f
C1010 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__conb_1_30/HI 3.81e-20
C1011 transmission_gate_9/GN V_HIGH 25.5f
C1012 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__inv_1_33/Y 0.0109f
C1013 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# 1.71e-19
C1014 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__inv_1_2/Y 0.0244f
C1015 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 5.18e-19
C1016 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_33/Y 3.89e-19
C1017 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 7.72e-20
C1018 sky130_fd_sc_hd__dfbbn_1_31/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0154f
C1019 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 6.71e-19
C1020 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 4.56e-21
C1021 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00141f
C1022 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# -2.65e-20
C1023 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.52e-19
C1024 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 8.14e-20
C1025 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.0291f
C1026 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 4.21e-21
C1027 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 1.87e-22
C1028 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__inv_1_9/Y 0.016f
C1029 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_21/Y 5.49e-20
C1030 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0111f
C1031 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# V_LOW 0.00802f
C1032 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q -1.38e-20
C1033 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 2.02e-20
C1034 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.6e-20
C1035 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_67/A 0.104f
C1036 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 3.84e-20
C1037 RISING_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 8.03e-21
C1038 sky130_fd_sc_hd__inv_1_36/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.267f
C1039 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.00155f
C1040 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0199f
C1041 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__nand2_8_9/A 1.7e-19
C1042 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.73e-19
C1043 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 1.48e-20
C1044 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.00208f
C1045 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_581_47# -2.6e-20
C1046 sky130_fd_sc_hd__dfbbn_1_21/Q_N FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.72e-19
C1047 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# V_LOW 0.0201f
C1048 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__inv_1_28/Y 0.0174f
C1049 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_1_49/Y 3.68e-21
C1050 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 7.5e-19
C1051 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 3.45e-20
C1052 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_193_47# 9.22e-20
C1053 Reset sky130_fd_sc_hd__inv_1_48/Y 0.205f
C1054 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 0.00369f
C1055 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_48/Y 0.0274f
C1056 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__inv_1_69/Y 1.05e-20
C1057 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__conb_1_37/HI 7.82e-19
C1058 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 6.53e-20
C1059 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 6.03e-20
C1060 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1_50/HI 2.62e-19
C1061 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# 0.00178f
C1062 sky130_fd_sc_hd__inv_1_3/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0173f
C1063 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__inv_1_36/Y 4.43e-21
C1064 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 5.11e-19
C1065 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0.0379f
C1066 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 5.35e-20
C1067 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# -1.24e-20
C1068 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.44e-21
C1069 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 7.65e-21
C1070 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 2.45e-20
C1071 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0294f
C1072 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1_45/LO 2.54e-21
C1073 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.111f
C1074 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_1_36/Y 1.37e-21
C1075 sky130_fd_sc_hd__inv_16_29/Y V_LOW 0.364f
C1076 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# V_LOW 0.00492f
C1077 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.028f
C1078 FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.15e-20
C1079 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 2.33e-19
C1080 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# sky130_fd_sc_hd__inv_16_41/Y 4.82e-20
C1081 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0258f
C1082 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_1_10/Y 0.0158f
C1083 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# -0.00385f
C1084 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__conb_1_47/HI 4.25e-19
C1085 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__inv_1_59/Y 0.00202f
C1086 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# V_LOW 2.94e-20
C1087 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_20/Y 0.048f
C1088 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# -6.23e-21
C1089 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -6.22e-19
C1090 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# -0.00463f
C1091 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1_34/LO 2.45e-21
C1092 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# Reset 0.00421f
C1093 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__inv_1_44/A 9.31e-19
C1094 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_581_47# 2.02e-19
C1095 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.0706f
C1096 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# V_LOW 4.8e-20
C1097 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_1_36/Y 4.74e-20
C1098 sky130_fd_sc_hd__inv_1_66/A Reset 0.0028f
C1099 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_27/Y 4e-20
C1100 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# V_LOW 0.00722f
C1101 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__nand2_1_5/Y 3.7e-20
C1102 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 9.33e-19
C1103 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/Q_N 1.16e-21
C1104 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00112f
C1105 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__nor2_1_0/Y 3.87e-20
C1106 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.127f
C1107 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00867f
C1108 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# -0.00782f
C1109 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0.027f
C1110 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 6.21e-20
C1111 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 2.93e-20
C1112 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 0.00124f
C1113 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 9.44e-20
C1114 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__inv_1_26/Y 0.00309f
C1115 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__conb_1_34/HI 8.17e-20
C1116 sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_28/Y 0.00439f
C1117 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_1_67/A 4.56e-21
C1118 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 0.00125f
C1119 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 2.09e-20
C1120 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 9.44e-19
C1121 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# sky130_fd_sc_hd__inv_16_40/Y 0.00181f
C1122 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_37/HI 2.75e-19
C1123 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 1.69e-19
C1124 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_24/Y 6.92e-19
C1125 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00294f
C1126 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_20/LO 5e-20
C1127 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# -3.86e-20
C1128 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# -0.0074f
C1129 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00162f
C1130 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# V_LOW 2.94e-20
C1131 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_30/HI 0.0108f
C1132 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 6.71e-19
C1133 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.03e-19
C1134 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__inv_1_12/Y 6.02e-19
C1135 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.36e-20
C1136 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_33/Y 6.56e-19
C1137 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_53/Y 0.0367f
C1138 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_21/HI 0.162f
C1139 sky130_fd_sc_hd__inv_16_22/A sky130_fd_sc_hd__inv_16_28/Y 1.35e-19
C1140 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# V_LOW 0.0217f
C1141 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.17e-19
C1142 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 0.00342f
C1143 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.00366f
C1144 sky130_fd_sc_hd__inv_1_49/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 2.5e-21
C1145 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.0103f
C1146 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_40/HI 0.001f
C1147 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 1.02e-20
C1148 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_52/A 4.01e-20
C1149 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.013f
C1150 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__inv_1_27/Y 4.95e-19
C1151 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.43e-21
C1152 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_19/Y 0.00857f
C1153 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# V_LOW -0.00169f
C1154 sky130_fd_sc_hd__dfbbn_1_18/a_581_47# sky130_fd_sc_hd__inv_1_28/Y 2.47e-19
C1155 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 7.72e-21
C1156 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_64/A 8.64e-20
C1157 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00147f
C1158 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00188f
C1159 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# 8.26e-21
C1160 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# V_LOW 0.0127f
C1161 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# 0.00159f
C1162 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__conb_1_3/HI 0.00351f
C1163 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.416f
C1164 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0224f
C1165 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.65e-20
C1166 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__conb_1_47/HI 1.05e-19
C1167 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 8.74e-19
C1168 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0187f
C1169 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 0.0711f
C1170 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__inv_1_30/Y 1.43e-21
C1171 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.66e-19
C1172 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_581_47# -2.6e-20
C1173 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# -6.43e-20
C1174 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# -3.06e-20
C1175 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 1.71e-21
C1176 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00143f
C1177 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_45/Y 0.0687f
C1178 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__inv_1_36/Y 2.52e-21
C1179 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0542f
C1180 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__nand2_8_1/a_27_47# 3.96e-19
C1181 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 1.91e-21
C1182 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_19/Y 0.342f
C1183 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__inv_1_35/Y 1.56e-20
C1184 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 3.13e-19
C1185 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# V_LOW 0.021f
C1186 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_22/Y 5.47e-19
C1187 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF17.Q 0.667f
C1188 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# -3.79e-20
C1189 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# -4.66e-20
C1190 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_1_43/Y 0.0211f
C1191 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_29/A 0.0197f
C1192 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_45/HI 0.049f
C1193 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_8/HI 0.0211f
C1194 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.62e-22
C1195 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 3.44e-20
C1196 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_16_40/Y 1.02e-19
C1197 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.25e-20
C1198 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_17/HI 6.95e-19
C1199 sky130_fd_sc_hd__conb_1_22/LO V_LOW 0.104f
C1200 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 7.54e-19
C1201 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.019f
C1202 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_581_47# -2.6e-20
C1203 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__conb_1_34/HI 0.0129f
C1204 sky130_fd_sc_hd__inv_16_55/Y CLOCK_GEN.SR_Op.Q 0.0635f
C1205 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_20/Y 4.97e-19
C1206 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/Q_N 1.17e-19
C1207 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nand2_1_5/Y 1.52e-19
C1208 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 1.34e-20
C1209 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_19/Y 3.16e-21
C1210 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1_67/A 1.63e-20
C1211 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_19/LO 8.84e-20
C1212 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_27_47# 2.03e-19
C1213 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0263f
C1214 sky130_fd_sc_hd__conb_1_11/LO V_LOW 0.133f
C1215 FALLING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 6.62f
C1216 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_3/HI 0.0119f
C1217 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0483f
C1218 sky130_fd_sc_hd__conb_1_26/LO FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00654f
C1219 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# -9.41e-19
C1220 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 4.49e-20
C1221 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_48/Y 0.00509f
C1222 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_2_0/A 3.62e-20
C1223 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__conb_1_19/HI -6.82e-19
C1224 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 5.26e-19
C1225 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 5.26e-19
C1226 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0164f
C1227 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__inv_1_12/Y 3.24e-19
C1228 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0123f
C1229 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF17.Q 0.317f
C1230 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__conb_1_21/HI -1.8e-19
C1231 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__conb_1_34/LO 1.38e-21
C1232 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# 7.83e-19
C1233 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# 8.4e-20
C1234 sky130_fd_sc_hd__inv_16_48/A sky130_fd_sc_hd__inv_16_50/A 2.16f
C1235 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.84e-19
C1236 sky130_fd_sc_hd__nor2_1_0/a_109_297# Reset 0.00167f
C1237 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.43e-19
C1238 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 2.01e-20
C1239 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 7.2e-19
C1240 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__conb_1_42/LO 9.17e-19
C1241 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 9.11e-19
C1242 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 0.026f
C1243 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_1_35/Y 8.09e-20
C1244 RISING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 1.89f
C1245 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.24e-19
C1246 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.23e-19
C1247 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# V_LOW 5.62e-20
C1248 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_1_22/Y 1.48e-20
C1249 sky130_fd_sc_hd__inv_1_56/A V_LOW 0.517f
C1250 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__inv_1_62/Y 6.69e-20
C1251 sky130_fd_sc_hd__dfbbn_1_1/Q_N FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00163f
C1252 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# -0.00336f
C1253 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# -3.79e-20
C1254 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# V_LOW -0.00121f
C1255 sky130_fd_sc_hd__conb_1_50/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 2.7e-19
C1256 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 7.73e-19
C1257 sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_44/A 0.00373f
C1258 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 0.0355f
C1259 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# sky130_fd_sc_hd__conb_1_47/HI 0.00138f
C1260 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 7.2e-19
C1261 FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.39f
C1262 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.21e-20
C1263 FALLING_COUNTER.COUNT_SUB_DFF6.Q V_LOW 1.93f
C1264 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__conb_1_25/HI 8.94e-20
C1265 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__inv_1_62/Y 3.47e-21
C1266 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 1.24e-19
C1267 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.12e-20
C1268 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.99e-19
C1269 CLOCK_GEN.SR_Op.Q FULL_COUNTER.COUNT_SUB_DFF0.Q 1.46e-20
C1270 sky130_fd_sc_hd__dfbbn_1_44/Q_N V_LOW -0.00509f
C1271 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 2.31e-19
C1272 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_25/Y 5.22e-20
C1273 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 0.369f
C1274 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# V_LOW 0.00462f
C1275 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# V_LOW 0.00883f
C1276 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -4.98e-19
C1277 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# -0.0103f
C1278 sky130_fd_sc_hd__conb_1_27/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0222f
C1279 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_26/Y 0.00224f
C1280 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# sky130_fd_sc_hd__inv_1_41/Y 7.97e-21
C1281 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF17.Q 3.93e-20
C1282 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_58/Y 0.207f
C1283 sky130_fd_sc_hd__conb_1_47/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0481f
C1284 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__conb_1_23/HI 7.9e-20
C1285 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__inv_1_31/Y 0.0771f
C1286 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_16_19/Y 0.00191f
C1287 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# -0.0103f
C1288 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# -0.00224f
C1289 sky130_fd_sc_hd__conb_1_34/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.71e-19
C1290 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_50/A 0.265f
C1291 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_66/A 3.04e-19
C1292 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__conb_1_35/HI 2.94e-20
C1293 sky130_fd_sc_hd__conb_1_12/HI FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0799f
C1294 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__nand2_1_5/Y 0.0287f
C1295 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__conb_1_17/HI 3.6e-21
C1296 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__conb_1_38/HI 0.00235f
C1297 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0287f
C1298 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_25/Y 0.0699f
C1299 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00887f
C1300 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_27/HI -0.00115f
C1301 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__conb_1_20/HI 7.4e-20
C1302 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# 0.00142f
C1303 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_0/HI 0.0407f
C1304 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__conb_1_9/HI 6.08e-20
C1305 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_381_47# -0.00516f
C1306 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__conb_1_37/HI 0.0113f
C1307 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.38e-19
C1308 RISING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0298f
C1309 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00309f
C1310 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# -0.00263f
C1311 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# -5.54e-21
C1312 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0141f
C1313 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__conb_1_19/HI -1.25e-20
C1314 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_27/Y 0.00307f
C1315 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__inv_1_34/Y 0.0108f
C1316 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 3.22e-20
C1317 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_791_47# 3.22e-20
C1318 sky130_fd_sc_hd__inv_16_44/Y CLOCK_GEN.SR_Op.Q 0.0616f
C1319 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 5.82e-19
C1320 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.00123f
C1321 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 1.53e-19
C1322 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 1.68e-19
C1323 RISING_COUNTER.COUNT_SUB_DFF12.Q V_LOW 2.17f
C1324 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.00157f
C1325 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.9e-20
C1326 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.00489f
C1327 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# V_LOW 0.0254f
C1328 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_50/A 0.158f
C1329 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__conb_1_21/HI -0.0089f
C1330 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 5.29e-19
C1331 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_31/Y 7.4e-19
C1332 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 5.57e-20
C1333 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 0.179f
C1334 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0.00837f
C1335 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# sky130_fd_sc_hd__conb_1_24/HI 8.26e-19
C1336 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__inv_1_38/Y 9.69e-19
C1337 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_1_64/A 0.00138f
C1338 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# Reset 0.00122f
C1339 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__nand2_8_4/Y 0.00154f
C1340 sky130_fd_sc_hd__dfbbn_1_2/Q_N V_LOW -0.00509f
C1341 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__inv_1_22/Y 8.92e-20
C1342 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__conb_1_30/HI 6.8e-21
C1343 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_891_329# 1.36e-21
C1344 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# V_LOW 0.0135f
C1345 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 6.53e-20
C1346 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 6.03e-20
C1347 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# sky130_fd_sc_hd__inv_1_48/Y 1.65e-21
C1348 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_12/LO 6.75e-21
C1349 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.132f
C1350 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_19/Y 0.00407f
C1351 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# 2.78e-21
C1352 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00133f
C1353 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 8.52e-19
C1354 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.43e-19
C1355 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF15.Q 0.02f
C1356 sky130_fd_sc_hd__inv_1_36/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0365f
C1357 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__inv_1_35/Y 2.81e-21
C1358 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 2.77e-20
C1359 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_68/Y 0.0043f
C1360 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# -6.8e-19
C1361 sky130_fd_sc_hd__inv_1_24/Y CLOCK_GEN.SR_Op.Q 0.0019f
C1362 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 5.58e-20
C1363 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 2.2e-20
C1364 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 4.49e-20
C1365 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 3.26e-19
C1366 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 1.98e-19
C1367 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00545f
C1368 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.00138f
C1369 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 9.2e-20
C1370 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0.00378f
C1371 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_48/Y 2.37e-19
C1372 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_3/A 9.63e-19
C1373 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nor2_1_0/Y 2.37e-20
C1374 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_557_413# -3.67e-20
C1375 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# -6.29e-19
C1376 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_2_0/A 6.31e-20
C1377 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# -9.41e-19
C1378 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_61/Y 0.376f
C1379 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 0.08f
C1380 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_193_47# 0.0301f
C1381 sky130_fd_sc_hd__conb_1_45/HI RISING_COUNTER.COUNT_SUB_DFF10.Q -4.84e-36
C1382 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0.0127f
C1383 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# V_LOW 4.8e-20
C1384 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.899f
C1385 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.93e-21
C1386 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__conb_1_17/HI 2.55e-19
C1387 sky130_fd_sc_hd__inv_16_15/Y sky130_fd_sc_hd__inv_16_32/Y 0.0403f
C1388 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 8.25e-19
C1389 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# 4.44e-19
C1390 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 5.34e-19
C1391 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_27/HI -2.07e-19
C1392 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__conb_1_20/HI 1.69e-19
C1393 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# V_LOW 0.0661f
C1394 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# 3.45e-20
C1395 sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0637f
C1396 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# V_LOW 2.26e-20
C1397 sky130_fd_sc_hd__conb_1_29/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 0.166f
C1398 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# -0.00107f
C1399 sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0309f
C1400 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# -0.00117f
C1401 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# -0.00149f
C1402 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# -9.32e-20
C1403 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0255f
C1404 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__nor2_1_0/Y 5.5e-21
C1405 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.022f
C1406 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# -8.61e-20
C1407 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.29e-20
C1408 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_791_47# 1.78e-20
C1409 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 1.78e-20
C1410 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 0.0228f
C1411 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# 2.32e-19
C1412 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0433f
C1413 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__inv_16_40/Y 2.86e-19
C1414 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_1_26/Y 0.00172f
C1415 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_1_49/Y 0.0105f
C1416 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 4.19e-20
C1417 sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_64/Y 1.28e-19
C1418 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# V_LOW -0.323f
C1419 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# V_LOW 2.94e-20
C1420 sky130_fd_sc_hd__inv_16_7/Y V_LOW 0.22f
C1421 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 1.95e-21
C1422 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00231f
C1423 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.67e-19
C1424 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_64/A 1.69e-20
C1425 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.78e-19
C1426 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__conb_1_51/HI 2.83e-20
C1427 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00338f
C1428 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 4.4e-19
C1429 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__conb_1_12/HI -0.0071f
C1430 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_37/Y 0.0254f
C1431 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 2.36e-20
C1432 FULL_COUNTER.COUNT_SUB_DFF6.Q V_LOW 3.94f
C1433 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.0243f
C1434 sky130_fd_sc_hd__dfbbn_1_9/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 5.89e-19
C1435 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 1.14e-19
C1436 sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF15.Q 8.52e-20
C1437 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# -2.37e-19
C1438 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# -3.88e-19
C1439 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_24/A 2.3e-19
C1440 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_8_4/Y 0.0222f
C1441 sky130_fd_sc_hd__nand2_8_2/a_27_47# Reset 0.1f
C1442 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__conb_1_10/HI 0.0207f
C1443 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 6.74e-20
C1444 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 8.67e-19
C1445 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 0.00384f
C1446 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 4.17e-20
C1447 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.00136f
C1448 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__conb_1_29/HI 0.0118f
C1449 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__conb_1_9/LO 8.31e-20
C1450 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0335f
C1451 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 2.87e-20
C1452 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 8.56e-21
C1453 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__conb_1_26/HI 2.17e-19
C1454 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 3.46e-21
C1455 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00198f
C1456 sky130_fd_sc_hd__conb_1_41/LO FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.89e-21
C1457 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_15/Y 0.16f
C1458 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_64/A 7.18e-20
C1459 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__inv_1_33/Y 9.49e-19
C1460 V_SENSE sky130_fd_sc_hd__conb_1_40/LO 9.19e-19
C1461 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI 0.00385f
C1462 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.00168f
C1463 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__conb_1_43/HI 0.0201f
C1464 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# Reset 6.6e-19
C1465 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__conb_1_25/LO 5.58e-20
C1466 sky130_fd_sc_hd__inv_1_55/Y V_LOW 0.154f
C1467 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_891_329# -2.2e-20
C1468 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# -0.00482f
C1469 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__nand3_1_2/Y 1.27e-19
C1470 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00629f
C1471 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# -0.01f
C1472 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_557_413# -3.67e-20
C1473 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# sky130_fd_sc_hd__conb_1_4/HI -6.57e-19
C1474 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 7.53e-20
C1475 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.00755f
C1476 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_47/Y 0.016f
C1477 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.114f
C1478 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 1.38e-20
C1479 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# 2e-19
C1480 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_381_47# -0.00516f
C1481 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_193_47# 3.1e-21
C1482 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.74e-20
C1483 sky130_fd_sc_hd__inv_16_42/Y Reset 0.0444f
C1484 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_66/Y 0.00211f
C1485 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_791_47# 0.00222f
C1486 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 1.86e-21
C1487 sky130_fd_sc_hd__conb_1_43/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.58e-19
C1488 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 6.67e-20
C1489 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.0223f
C1490 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_18/A 1.78e-20
C1491 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__conb_1_20/HI 0.00116f
C1492 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_23/HI 2.49e-21
C1493 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# -3.8e-20
C1494 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# -5.54e-21
C1495 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# V_LOW 0.00546f
C1496 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 8.84e-20
C1497 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# V_LOW 2.94e-20
C1498 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__conb_1_46/HI -0.0016f
C1499 sky130_fd_sc_hd__inv_1_67/A V_LOW 1.13f
C1500 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# V_LOW 0.0114f
C1501 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_8_0/Y 0.0015f
C1502 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.137f
C1503 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__conb_1_5/HI 2.38e-19
C1504 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 3.34e-19
C1505 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_1_12/Y 3.61e-21
C1506 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/Q_N -4.78e-20
C1507 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_23/HI 0.00145f
C1508 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_55/A 1.07f
C1509 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 4.31e-23
C1510 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__inv_1_32/Y 0.00209f
C1511 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 8.17e-20
C1512 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_581_47# -7.91e-19
C1513 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00123f
C1514 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.81e-20
C1515 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# V_LOW 0.00635f
C1516 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__conb_1_11/HI 4.72e-19
C1517 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__conb_1_45/HI 1.03e-19
C1518 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.582f
C1519 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.22e-19
C1520 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# sky130_fd_sc_hd__inv_1_26/Y 5.8e-19
C1521 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.45e-20
C1522 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 2.44e-20
C1523 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 1.35e-20
C1524 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 1.44e-20
C1525 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_557_413# 1e-19
C1526 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0342f
C1527 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__conb_1_12/HI 8.88e-20
C1528 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.06e-19
C1529 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 6.36e-20
C1530 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__inv_1_38/Y 2.22e-20
C1531 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__nand2_8_8/A 0.00371f
C1532 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 9.23e-19
C1533 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_30/HI 0.08f
C1534 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_473_413# -4.53e-19
C1535 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 4.88e-21
C1536 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__conb_1_32/HI -0.048f
C1537 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# V_LOW 0.0126f
C1538 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# -1.66e-19
C1539 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.003f
C1540 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 9.05e-19
C1541 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 8.4e-21
C1542 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 6.66e-19
C1543 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# -0.0395f
C1544 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# sky130_fd_sc_hd__conb_1_10/HI 4.96e-20
C1545 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 3.78e-19
C1546 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__conb_1_29/HI 0.0203f
C1547 RISING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.2f
C1548 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__conb_1_26/HI 5.26e-19
C1549 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 0.021f
C1550 FULL_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.027f
C1551 sky130_fd_sc_hd__inv_1_32/Y FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.47e-19
C1552 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__conb_1_50/HI 0.0218f
C1553 sky130_fd_sc_hd__dfbbn_1_46/a_557_413# sky130_fd_sc_hd__inv_1_50/Y 8.17e-19
C1554 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 3.19e-19
C1555 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# -0.00869f
C1556 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand3_1_2/Y 0.00765f
C1557 sky130_fd_sc_hd__conb_1_5/LO V_LOW 0.187f
C1558 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__conb_1_44/HI 4.93e-19
C1559 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__inv_1_41/Y 0.044f
C1560 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__conb_1_29/HI 6.93e-21
C1561 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__conb_1_43/HI 2.47e-21
C1562 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00907f
C1563 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# -3.46e-20
C1564 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# -4.33e-19
C1565 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 2.66e-19
C1566 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 5.75e-19
C1567 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/Q_N 2.89e-19
C1568 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0104f
C1569 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00252f
C1570 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__conb_1_23/HI 5.13e-20
C1571 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# -0.00107f
C1572 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 1.21e-20
C1573 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 3.97e-22
C1574 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 4.23e-20
C1575 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 3.16e-21
C1576 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00861f
C1577 sky130_fd_sc_hd__dfbbn_1_0/Q_N FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00231f
C1578 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.45e-21
C1579 sky130_fd_sc_hd__inv_1_7/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0148f
C1580 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.041f
C1581 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 0.0224f
C1582 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.128f
C1583 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_891_329# -2.2e-20
C1584 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -4.72e-19
C1585 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.05e-19
C1586 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 0.0354f
C1587 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# -9.32e-20
C1588 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 9.37e-21
C1589 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_941_21# -1.62e-20
C1590 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# -2.32e-19
C1591 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 5.48e-21
C1592 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_47/Y 2.68e-21
C1593 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF14.Q 0.369f
C1594 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0379f
C1595 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_4/Y 5.64e-21
C1596 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__inv_1_40/Y 1.02e-20
C1597 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_19/LO 0.0223f
C1598 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_22/Y 8.12e-22
C1599 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 0.0224f
C1600 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_28/HI 0.0315f
C1601 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_381_47# -2.53e-20
C1602 sky130_fd_sc_hd__nand2_1_3/Y CLOCK_GEN.SR_Op.Q 7.73e-20
C1603 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_44/A 2.66e-19
C1604 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_33/LO 2.01e-20
C1605 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__conb_1_45/HI 1.65e-20
C1606 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 4.55e-20
C1607 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_1_5/Y 0.0528f
C1608 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__inv_1_49/Y 1.31e-22
C1609 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__conb_1_32/HI 0.03f
C1610 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__conb_1_5/HI -0.00233f
C1611 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 2.41e-19
C1612 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.00893f
C1613 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_33/Y 5.08e-21
C1614 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 3.86e-20
C1615 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_52/A 2.88e-21
C1616 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 9.36e-21
C1617 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_31/HI 0.00546f
C1618 sky130_fd_sc_hd__inv_1_45/Y V_LOW 0.466f
C1619 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.79e-20
C1620 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__inv_16_40/Y 0.114f
C1621 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__conb_1_19/HI 1.11e-19
C1622 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 7.46e-21
C1623 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 8.3e-19
C1624 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_25/LO 0.00869f
C1625 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# sky130_fd_sc_hd__inv_1_44/A 2.83e-19
C1626 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__conb_1_12/HI -1.27e-19
C1627 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 4.16e-19
C1628 sky130_fd_sc_hd__conb_1_12/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 0.024f
C1629 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_47/Y 0.001f
C1630 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# -0.00116f
C1631 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 0.0633f
C1632 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 0.00184f
C1633 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__conb_1_8/HI 1.1e-22
C1634 sky130_fd_sc_hd__conb_1_26/LO FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.57e-20
C1635 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__conb_1_29/HI 0.0278f
C1636 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_1_13/Y 8.36e-19
C1637 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0.00421f
C1638 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# 3.77e-19
C1639 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00874f
C1640 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00291f
C1641 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__conb_1_26/HI 9.57e-19
C1642 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__inv_1_12/Y 1.67e-19
C1643 sky130_fd_sc_hd__inv_1_25/Y sky130_fd_sc_hd__inv_1_28/Y 2.11e-19
C1644 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__conb_1_21/HI 6.34e-21
C1645 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# V_LOW 5.11e-19
C1646 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# -0.00141f
C1647 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__inv_1_10/Y 4.29e-20
C1648 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# V_LOW 2.26e-20
C1649 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00252f
C1650 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_1_45/Y 0.00122f
C1651 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_56/A 1.77e-21
C1652 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__inv_1_29/Y 4.75e-20
C1653 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.63e-19
C1654 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.266f
C1655 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# V_LOW -9.15e-19
C1656 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.3e-19
C1657 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 0.00625f
C1658 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 5.66e-20
C1659 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0302f
C1660 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.26f
C1661 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_64/Y 0.00215f
C1662 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# V_LOW 0.0194f
C1663 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_2_0/A 0.00404f
C1664 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# V_LOW 0.0081f
C1665 sky130_fd_sc_hd__inv_1_20/Y V_LOW 0.179f
C1666 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/Q_N 2.55e-21
C1667 sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 0.00128f
C1668 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00707f
C1669 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_8/HI 9.3e-19
C1670 sky130_fd_sc_hd__inv_16_2/Y Reset 0.0561f
C1671 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# -0.00471f
C1672 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# -0.00336f
C1673 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# -3.79e-20
C1674 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 1.87e-20
C1675 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_1_69/Y 1.72e-20
C1676 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__inv_1_8/Y 3.92e-20
C1677 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_9/HI 0.0307f
C1678 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__conb_1_38/LO 4.39e-20
C1679 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/Q_N -4.78e-20
C1680 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0085f
C1681 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# -1.66e-19
C1682 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_791_47# -2.22e-34
C1683 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 8.26e-21
C1684 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__conb_1_32/HI 6.34e-20
C1685 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0461f
C1686 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_66/A 0.0247f
C1687 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# V_LOW 1.38e-19
C1688 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_2/Y 0.136f
C1689 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.00264f
C1690 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_42/Y 0.0864f
C1691 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF14.Q 0.276f
C1692 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_193_47# -0.0586f
C1693 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# -0.00141f
C1694 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 5.48e-21
C1695 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__nand2_1_2/A 1.14e-20
C1696 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__inv_1_25/Y 6.73e-20
C1697 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1_16/HI 0.0225f
C1698 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 0.106f
C1699 sky130_fd_sc_hd__conb_1_33/HI V_LOW 0.0287f
C1700 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_19/LO 6.66e-19
C1701 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# sky130_fd_sc_hd__conb_1_32/HI 5.18e-19
C1702 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# sky130_fd_sc_hd__conb_1_5/HI -0.00261f
C1703 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__inv_1_61/Y 0.00477f
C1704 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 1.49e-19
C1705 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 8.12e-19
C1706 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 7.19e-19
C1707 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 9.78e-19
C1708 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0202f
C1709 sky130_fd_sc_hd__inv_16_6/A FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0309f
C1710 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# Reset 0.0562f
C1711 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.04e-21
C1712 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# sky130_fd_sc_hd__conb_1_19/HI 1.66e-20
C1713 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__conb_1_25/LO 0.00169f
C1714 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__conb_1_23/HI -0.00175f
C1715 sky130_fd_sc_hd__conb_1_45/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00852f
C1716 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0.0403f
C1717 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# -3.69e-19
C1718 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# -0.00139f
C1719 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# -0.00985f
C1720 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# -0.00631f
C1721 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__conb_1_3/HI 2.76e-19
C1722 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__conb_1_10/HI 1.18e-20
C1723 V_SENSE sky130_fd_sc_hd__conb_1_40/HI 6.59e-19
C1724 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI 0.0242f
C1725 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 9.95e-20
C1726 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 5.19e-19
C1727 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0634f
C1728 sky130_fd_sc_hd__inv_1_3/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0268f
C1729 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 0.00104f
C1730 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_8/LO 9.67e-19
C1731 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00609f
C1732 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__inv_1_31/Y 0.00102f
C1733 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 2.92e-19
C1734 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 1.03e-19
C1735 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00251f
C1736 sky130_fd_sc_hd__dfbbn_1_47/a_581_47# sky130_fd_sc_hd__inv_1_45/Y 5.8e-19
C1737 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.19e-20
C1738 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_49/Y 0.0727f
C1739 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 4.07e-19
C1740 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__conb_1_11/HI 0.00592f
C1741 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_59/Y 0.0765f
C1742 sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16_49/A 0.0955f
C1743 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 1.1e-19
C1744 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 6.32e-19
C1745 sky130_fd_sc_hd__conb_1_22/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0231f
C1746 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 8.17e-19
C1747 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0074f
C1748 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_56/Y 0.125f
C1749 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/Q_N 1.31e-19
C1750 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__inv_1_10/Y 0.0417f
C1751 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__conb_1_27/HI 3.51e-20
C1752 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_64/Y 2.31e-19
C1753 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# V_LOW 2.94e-20
C1754 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_381_47# -3.03e-19
C1755 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# -6.23e-21
C1756 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_891_329# 0.00181f
C1757 sky130_fd_sc_hd__dfbbn_1_40/Q_N FALLING_COUNTER.COUNT_SUB_DFF7.Q 6.87e-19
C1758 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# sky130_fd_sc_hd__conb_1_33/HI -6.57e-19
C1759 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_2_0/A 0.102f
C1760 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__conb_1_7/HI 4.32e-21
C1761 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_16_40/Y 0.00111f
C1762 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0754f
C1763 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 6.6e-20
C1764 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__conb_1_23/HI 0.0152f
C1765 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0399f
C1766 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.76e-20
C1767 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 3.33e-20
C1768 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__inv_1_40/Y 2.2e-19
C1769 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# 1.4e-19
C1770 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_8_9/A 0.00424f
C1771 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_34/LO 0.0283f
C1772 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00802f
C1773 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 8.26e-21
C1774 sky130_fd_sc_hd__dfbbn_1_45/Q_N RISING_COUNTER.COUNT_SUB_DFF4.Q 5.1e-20
C1775 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 2.02e-21
C1776 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 9.02e-19
C1777 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 3.3e-19
C1778 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 2.16e-19
C1779 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__conb_1_2/HI 0.00243f
C1780 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# V_LOW 0.0171f
C1781 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_32/HI 0.00195f
C1782 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 8.56e-20
C1783 sky130_fd_sc_hd__conb_1_22/HI FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00203f
C1784 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0998f
C1785 V_SENSE sky130_fd_sc_hd__inv_16_55/A 0.00544f
C1786 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 5.01e-19
C1787 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 1.98e-20
C1788 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# V_LOW 1.38e-19
C1789 sky130_fd_sc_hd__inv_16_20/A sky130_fd_sc_hd__inv_16_19/Y 4.33e-20
C1790 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# Reset 3.47e-19
C1791 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0649f
C1792 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# V_LOW 3.96e-19
C1793 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_38/HI 0.00401f
C1794 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__inv_1_1/Y 0.00318f
C1795 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_791_47# 2.22e-34
C1796 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# -1.76e-19
C1797 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0677f
C1798 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.18e-19
C1799 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 5.1e-19
C1800 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__conb_1_3/HI 7.03e-19
C1801 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_23/HI 0.00263f
C1802 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__inv_1_60/Y 2.47e-20
C1803 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_30/HI 0.00215f
C1804 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# -6.43e-20
C1805 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# -3.06e-20
C1806 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 2.2e-20
C1807 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.00968f
C1808 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.0396f
C1809 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_1_13/Y 0.0107f
C1810 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.152f
C1811 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# V_LOW 0.0131f
C1812 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__inv_1_14/Y 1.07e-20
C1813 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_16_40/Y 0.0451f
C1814 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.601f
C1815 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# sky130_fd_sc_hd__conb_1_45/HI 2.43e-19
C1816 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__conb_1_41/HI -4.95e-19
C1817 sky130_fd_sc_hd__dfbbn_1_21/Q_N FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0137f
C1818 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00152f
C1819 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 6.82e-21
C1820 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_4/HI 0.0987f
C1821 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__conb_1_11/HI 0.0101f
C1822 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__inv_1_38/Y 0.0292f
C1823 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_45/Y 2.36e-21
C1824 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.66e-19
C1825 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_19/HI 6.75e-19
C1826 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0241f
C1827 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# sky130_fd_sc_hd__inv_1_10/Y 0.00117f
C1828 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# -1.69e-19
C1829 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 3.27e-19
C1830 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00137f
C1831 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 2.53e-19
C1832 sky130_fd_sc_hd__conb_1_44/LO FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00299f
C1833 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_53/A 0.004f
C1834 sky130_fd_sc_hd__dfbbn_1_12/Q_N V_LOW 1.99e-19
C1835 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__conb_1_47/HI 0.00457f
C1836 V_SENSE sky130_fd_sc_hd__inv_16_8/Y 0.0536f
C1837 sky130_fd_sc_hd__dfbbn_1_19/a_557_413# sky130_fd_sc_hd__inv_1_28/Y 8.17e-19
C1838 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_8_0/A 0.0254f
C1839 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_19/LO 3.11e-19
C1840 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# sky130_fd_sc_hd__inv_2_0/A 0.00147f
C1841 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 2.18e-19
C1842 sky130_fd_sc_hd__inv_16_6/A RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0308f
C1843 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.0597f
C1844 FULL_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.01f
C1845 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF8.Q 1.94e-20
C1846 RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 1.09f
C1847 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# -0.00125f
C1848 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# -0.00393f
C1849 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_12/HI 6.23e-20
C1850 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.96e-20
C1851 sky130_fd_sc_hd__nand2_1_2/A FULL_COUNTER.COUNT_SUB_DFF2.Q 4.48e-20
C1852 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_48/LO 9.65e-21
C1853 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00229f
C1854 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -0.0114f
C1855 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# -7.77e-19
C1856 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 2.63e-21
C1857 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.05e-19
C1858 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 3.3e-21
C1859 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 3.72e-21
C1860 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 1.61e-20
C1861 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__inv_1_55/Y 0.0375f
C1862 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__inv_16_40/Y 0.00157f
C1863 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.00509f
C1864 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 1.86e-21
C1865 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 6.59e-21
C1866 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00337f
C1867 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# sky130_fd_sc_hd__conb_1_2/HI 1.69e-19
C1868 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_66/Y 2.07e-20
C1869 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_25/LO 4.49e-20
C1870 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.00746f
C1871 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 6.31e-21
C1872 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.23e-21
C1873 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# V_LOW 0.00471f
C1874 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 2.27e-20
C1875 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_47/A 5.63e-19
C1876 sky130_fd_sc_hd__inv_1_7/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.524f
C1877 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# V_LOW 2.94e-20
C1878 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__conb_1_39/HI 1.07e-20
C1879 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# -6.43e-20
C1880 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# CLOCK_GEN.SR_Op.Q 0.00471f
C1881 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# -0.00985f
C1882 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_23/HI 0.0967f
C1883 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0309f
C1884 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.26e-19
C1885 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# V_LOW -0.00448f
C1886 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__inv_1_1/Y 1.07e-21
C1887 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_30/Y 0.069f
C1888 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 5.46e-20
C1889 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00132f
C1890 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 3.31e-19
C1891 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__inv_16_41/Y 0.0013f
C1892 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00147f
C1893 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 2.73e-20
C1894 sky130_fd_sc_hd__conb_1_39/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 8.4e-19
C1895 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0382f
C1896 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__conb_1_9/HI 3.09e-19
C1897 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 9.83e-21
C1898 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0283f
C1899 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.0351f
C1900 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 0.811f
C1901 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# V_LOW 4.77e-19
C1902 sky130_fd_sc_hd__conb_1_37/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0346f
C1903 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__inv_1_8/Y 1.31e-20
C1904 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__conb_1_12/HI 1.19e-19
C1905 sky130_fd_sc_hd__conb_1_45/HI sky130_fd_sc_hd__dfbbn_1_49/Q_N -2.17e-19
C1906 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_56/Y 0.0155f
C1907 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 0.00532f
C1908 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 4.27e-21
C1909 sky130_fd_sc_hd__conb_1_27/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0031f
C1910 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# sky130_fd_sc_hd__conb_1_4/HI 8.44e-20
C1911 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 3.01e-19
C1912 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# sky130_fd_sc_hd__inv_1_38/Y 5.29e-19
C1913 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__conb_1_51/HI 0.126f
C1914 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_62/Y 0.169f
C1915 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00269f
C1916 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0015f
C1917 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_581_47# -7.91e-19
C1918 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00837f
C1919 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__inv_1_32/Y 0.00112f
C1920 sky130_fd_sc_hd__inv_1_18/A V_LOW 0.397f
C1921 sky130_fd_sc_hd__conb_1_38/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00156f
C1922 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0358f
C1923 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0493f
C1924 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__conb_1_51/HI 2.38e-19
C1925 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.96e-19
C1926 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__conb_1_15/LO 1.85e-21
C1927 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_43/HI 0.508f
C1928 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__conb_1_44/HI 1.36e-20
C1929 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__inv_1_27/Y 0.0119f
C1930 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 5.81e-20
C1931 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# -2.52e-19
C1932 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -1.89e-19
C1933 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_2_0/A 1.17e-19
C1934 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 1.38e-19
C1935 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q -2.71e-20
C1936 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# sky130_fd_sc_hd__inv_1_44/A 3.56e-20
C1937 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 1.74e-20
C1938 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 1.61e-20
C1939 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__inv_1_35/Y 2.12e-19
C1940 sky130_fd_sc_hd__inv_16_40/Y transmission_gate_9/GN 5.03e-20
C1941 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# V_LOW -0.316f
C1942 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 0.0141f
C1943 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__conb_1_6/HI 5.68e-20
C1944 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 2e-19
C1945 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_48/Q_N 2.21e-20
C1946 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 7.65e-20
C1947 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 7.65e-20
C1948 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0031f
C1949 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# -1.66e-19
C1950 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00357f
C1951 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_1_0/a_113_47# 1.06e-19
C1952 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__inv_1_13/Y 0.172f
C1953 sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 4.48e-20
C1954 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0583f
C1955 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# sky130_fd_sc_hd__conb_1_15/HI 5.67e-19
C1956 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_23/Y 2.69e-19
C1957 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0.0171f
C1958 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__conb_1_2/HI 0.00926f
C1959 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_8/HI 0.00223f
C1960 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -6.22e-19
C1961 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# -6.23e-21
C1962 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# -0.00367f
C1963 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_16/HI 0.285f
C1964 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 2.3e-19
C1965 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# V_LOW 0.00924f
C1966 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0977f
C1967 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_1_26/Y 6.61e-19
C1968 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# V_LOW -0.114f
C1969 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_38/Q_N 4.68e-20
C1970 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.19e-20
C1971 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 8.17e-19
C1972 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# V_LOW 4.8e-20
C1973 V_SENSE sky130_fd_sc_hd__conb_1_41/LO 9.19e-19
C1974 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_30/Y 0.121f
C1975 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_1_29/Y 0.0367f
C1976 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 1.36e-19
C1977 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00152f
C1978 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.01e-20
C1979 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__conb_1_7/HI -0.00964f
C1980 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0421f
C1981 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# V_LOW 0.00567f
C1982 sky130_fd_sc_hd__conb_1_36/LO RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00196f
C1983 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__conb_1_20/HI -2.12e-19
C1984 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 0.0213f
C1985 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_51/Y 0.0028f
C1986 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1_45/LO 7.91e-19
C1987 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 0.0365f
C1988 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# V_LOW -0.00121f
C1989 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__conb_1_19/HI 8.54e-19
C1990 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_1_24/Y 5.83e-20
C1991 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__inv_1_14/Y 5.85e-22
C1992 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 8.06e-19
C1993 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_3/A 9.02e-19
C1994 sky130_fd_sc_hd__conb_1_32/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 1.91e-22
C1995 sky130_fd_sc_hd__conb_1_46/HI V_LOW 0.221f
C1996 sky130_fd_sc_hd__inv_1_36/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00343f
C1997 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_47/Y 2.59e-20
C1998 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/Y 0.00481f
C1999 sky130_fd_sc_hd__dfbbn_1_23/Q_N FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.68e-20
C2000 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 0.00114f
C2001 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_38/HI 0.0155f
C2002 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 0.0132f
C2003 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# V_LOW -0.118f
C2004 sky130_fd_sc_hd__inv_16_6/A FULL_COUNTER.COUNT_SUB_DFF1.Q 0.848f
C2005 sky130_fd_sc_hd__conb_1_16/HI sky130_fd_sc_hd__conb_1_15/HI 9.79e-20
C2006 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# V_LOW 4.8e-20
C2007 V_SENSE sky130_fd_sc_hd__fill_4_215/VPB 0.0446f
C2008 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0255f
C2009 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0209f
C2010 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.95e-19
C2011 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.324f
C2012 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__conb_1_51/HI 4.32e-20
C2013 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__inv_16_41/Y 5.28e-20
C2014 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0322f
C2015 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# V_LOW 0.0221f
C2016 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# 1.04e-19
C2017 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_791_47# -2.22e-34
C2018 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# -1.76e-19
C2019 sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 1.48e-19
C2020 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0311f
C2021 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 6.08e-20
C2022 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_5/HI 0.00339f
C2023 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.116f
C2024 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/Q_N -9.56e-20
C2025 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 0.00179f
C2026 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_17/HI 8.97e-19
C2027 sky130_fd_sc_hd__nand2_8_9/A V_LOW 0.0889f
C2028 sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# sky130_fd_sc_hd__conb_1_6/HI 0.00264f
C2029 FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0499f
C2030 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0212f
C2031 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_24/LO 0.0122f
C2032 sky130_fd_sc_hd__conb_1_39/LO RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0718f
C2033 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__conb_1_16/LO 8.81e-20
C2034 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_42/Y 0.277f
C2035 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0.0127f
C2036 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.9e-20
C2037 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 6.42e-20
C2038 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 4.5e-20
C2039 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 7.09e-19
C2040 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_22/LO 8.84e-20
C2041 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 0.0324f
C2042 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0011f
C2043 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_581_47# 3.08e-19
C2044 sky130_fd_sc_hd__nand3_1_1/Y V_LOW 0.231f
C2045 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_6/HI 1.21e-19
C2046 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 9.4e-19
C2047 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 4.17e-20
C2048 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 7.23e-20
C2049 V_SENSE sky130_fd_sc_hd__conb_1_43/LO 9.19e-19
C2050 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# -0.00441f
C2051 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 2.78e-21
C2052 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# V_LOW 0.00351f
C2053 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__conb_1_16/HI 0.00402f
C2054 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__inv_1_25/Y 6.14e-20
C2055 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# V_LOW -9.94e-19
C2056 sky130_fd_sc_hd__conb_1_6/HI V_LOW 0.124f
C2057 sky130_fd_sc_hd__dfbbn_1_9/Q_N FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00488f
C2058 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 0.00996f
C2059 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 3.58e-19
C2060 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# -0.0022f
C2061 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# -5.54e-21
C2062 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.381f
C2063 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__conb_1_7/HI -6.8e-19
C2064 sky130_fd_sc_hd__inv_1_67/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 1.46e-20
C2065 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 0.192f
C2066 sky130_fd_sc_hd__conb_1_3/HI FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0254f
C2067 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_64/A 5.54e-19
C2068 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.88e-20
C2069 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# sky130_fd_sc_hd__conb_1_20/HI -1.57e-20
C2070 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_581_47# 5.31e-19
C2071 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0295f
C2072 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.147f
C2073 sky130_fd_sc_hd__nand2_8_6/a_27_47# V_LOW -0.0117f
C2074 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00622f
C2075 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_16_4/Y 0.00382f
C2076 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 0.0034f
C2077 V_SENSE sky130_fd_sc_hd__inv_16_29/A 0.0241f
C2078 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# sky130_fd_sc_hd__inv_1_13/Y 1.88e-20
C2079 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 9.58e-21
C2080 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 2.85e-19
C2081 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__conb_1_50/HI 0.00506f
C2082 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# -2.53e-20
C2083 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0356f
C2084 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# 7.13e-19
C2085 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# -0.00889f
C2086 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 4.78e-20
C2087 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# V_LOW -9.94e-19
C2088 V_SENSE sky130_fd_sc_hd__inv_16_26/A 0.0535f
C2089 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 0.00519f
C2090 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__inv_16_41/Y 0.0227f
C2091 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_19/HI 0.00508f
C2092 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__inv_1_35/Y 0.0116f
C2093 sky130_fd_sc_hd__nand2_1_1/a_113_47# V_LOW -1.78e-19
C2094 sky130_fd_sc_hd__inv_16_55/A CLOCK_GEN.SR_Op.Q 0.0619f
C2095 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.11e-20
C2096 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.57e-19
C2097 sky130_fd_sc_hd__inv_8_0/A V_LOW 0.439f
C2098 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__conb_1_24/HI 7.32e-20
C2099 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# V_LOW -6.55e-19
C2100 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00245f
C2101 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00771f
C2102 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_53/A 0.0315f
C2103 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand3_1_2/a_193_47# 1.72e-19
C2104 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 9.99e-21
C2105 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 6.53e-19
C2106 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# 0.00211f
C2107 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_1_46/A 1.72e-19
C2108 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0408f
C2109 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_65/A 0.02f
C2110 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__nand2_1_2/A 3.24e-21
C2111 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.31e-19
C2112 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 9.48e-20
C2113 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 9.48e-20
C2114 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.21e-19
C2115 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.00352f
C2116 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 1.21e-19
C2117 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__conb_1_31/HI 1.61e-19
C2118 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_473_413# -0.00834f
C2119 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -5.02e-19
C2120 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 0.00895f
C2121 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_1_0/Y 0.00195f
C2122 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0711f
C2123 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__inv_16_40/Y 0.0246f
C2124 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# V_LOW -9.15e-19
C2125 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 9.32e-19
C2126 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# 7.22e-19
C2127 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# -0.00149f
C2128 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# -1.67e-19
C2129 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.168f
C2130 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 3.31e-20
C2131 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# -1.44e-20
C2132 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 4.68e-20
C2133 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 7.83e-20
C2134 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__conb_1_35/HI -0.00135f
C2135 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_40/HI -3.61e-19
C2136 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_473_413# 1.28e-19
C2137 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 7.41e-22
C2138 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 2.47e-21
C2139 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 7.25e-20
C2140 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__conb_1_46/HI 1.6e-19
C2141 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# V_LOW 0.0216f
C2142 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_8/HI 2.16e-20
C2143 V_SENSE sky130_fd_sc_hd__conb_1_45/HI 0.00156f
C2144 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# V_LOW 2.26e-20
C2145 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 4.58e-19
C2146 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 7.44e-21
C2147 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_791_47# 2.38e-20
C2148 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0277f
C2149 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# -0.0238f
C2150 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_557_413# -3.67e-20
C2151 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# -7.47e-20
C2152 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__conb_1_7/HI -2.17e-19
C2153 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 8.4e-21
C2154 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 6.66e-19
C2155 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.003f
C2156 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 9.05e-19
C2157 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0.0165f
C2158 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_25/HI 0.0294f
C2159 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_56/A 3.56e-19
C2160 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0.0375f
C2161 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 3.75e-20
C2162 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 3.75e-20
C2163 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.52e-19
C2164 RISING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.08f
C2165 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0646f
C2166 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_32/HI 3.38e-19
C2167 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_21/Y 1.17e-21
C2168 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_16/Y 1.12e-19
C2169 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 3.41e-19
C2170 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 5.61e-20
C2171 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 2.16e-19
C2172 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 2.35e-19
C2173 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 3.19e-21
C2174 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_23/HI 1.87e-21
C2175 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_1_26/Y 0.281f
C2176 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00778f
C2177 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_25/Y 0.13f
C2178 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__nor2_1_0/Y 0.3f
C2179 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 9.03e-21
C2180 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_15/HI 0.285f
C2181 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_16_40/Y 0.0026f
C2182 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.07e-20
C2183 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0331f
C2184 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__conb_1_27/HI 9.67e-20
C2185 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_193_47# -0.142f
C2186 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# V_LOW 1.38e-19
C2187 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_16_40/Y 0.0333f
C2188 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__conb_1_13/LO 1.22e-20
C2189 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# sky130_fd_sc_hd__conb_1_9/HI 2.4e-19
C2190 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_51/Y 1.04f
C2191 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# -0.00141f
C2192 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# 1.44e-21
C2193 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_64/A 1.53e-20
C2194 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.04f
C2195 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.25e-21
C2196 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_581_47# -2.6e-20
C2197 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.32f
C2198 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.8e-20
C2199 sky130_fd_sc_hd__inv_1_7/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 2.08e-19
C2200 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0242f
C2201 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0272f
C2202 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_33/Y 0.00605f
C2203 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00408f
C2204 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__conb_1_24/LO 0.00643f
C2205 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 0.00194f
C2206 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.04e-21
C2207 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__conb_1_14/HI 0.00205f
C2208 sky130_fd_sc_hd__inv_2_0/A V_LOW 2.4f
C2209 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_1_24/A 9.8e-19
C2210 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_63/Y 0.155f
C2211 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0216f
C2212 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 4.1e-19
C2213 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 1.2e-21
C2214 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 1.75e-21
C2215 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 9.2e-22
C2216 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 2.35e-20
C2217 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 8.72e-19
C2218 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00547f
C2219 sky130_fd_sc_hd__nand2_8_8/a_27_47# V_LOW -0.0117f
C2220 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__conb_1_39/HI -6.52e-20
C2221 sky130_fd_sc_hd__conb_1_37/HI FULL_COUNTER.COUNT_SUB_DFF0.Q 0.159f
C2222 Reset transmission_gate_9/GN 12.2f
C2223 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.75e-21
C2224 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_557_413# 5.03e-19
C2225 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__inv_1_50/Y 1.22e-20
C2226 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0416f
C2227 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_33/HI 1.88e-19
C2228 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# -0.00248f
C2229 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_16_2/Y 2.89e-19
C2230 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__conb_1_31/HI 2.12e-19
C2231 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# -2.57e-20
C2232 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_33/Y 6.77e-19
C2233 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 2.89e-20
C2234 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__inv_1_0/Y 9.37e-21
C2235 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.42e-19
C2236 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0569f
C2237 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__inv_1_14/Y 0.023f
C2238 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_46/A 0.1f
C2239 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# sky130_fd_sc_hd__inv_1_41/Y 0.00142f
C2240 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 2.55e-20
C2241 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__inv_1_59/Y 0.0574f
C2242 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# 1.06e-20
C2243 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI 2.08e-21
C2244 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 4.15e-20
C2245 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__conb_1_35/HI -2.07e-19
C2246 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__conb_1_40/HI 6.7e-21
C2247 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.53e-20
C2248 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.0151f
C2249 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.283f
C2250 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# -5.75e-19
C2251 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# -0.0103f
C2252 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -5.54e-21
C2253 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__inv_1_49/Y 0.00175f
C2254 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.14f
C2255 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_381_47# 2.27e-19
C2256 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.51e-19
C2257 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.1e-20
C2258 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/Q_N -4.78e-20
C2259 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 0.00507f
C2260 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00785f
C2261 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# -0.00774f
C2262 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_16_40/Y 7.09e-21
C2263 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 5.34e-19
C2264 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 5.34e-19
C2265 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.0601f
C2266 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 2.19e-20
C2267 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.16e-19
C2268 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_30/LO 5.04e-21
C2269 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 2.64e-19
C2270 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 0.00143f
C2271 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 7.14e-20
C2272 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 2.09e-19
C2273 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_791_47# 9.9e-20
C2274 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# sky130_fd_sc_hd__inv_1_26/Y 0.00252f
C2275 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_16_40/Y 3.45e-20
C2276 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 8.92e-21
C2277 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 0.02f
C2278 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# sky130_fd_sc_hd__inv_1_2/Y 3.75e-21
C2279 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# V_LOW 2.26e-20
C2280 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__conb_1_33/LO 9.82e-19
C2281 sky130_fd_sc_hd__conb_1_4/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0623f
C2282 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.00397f
C2283 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00591f
C2284 sky130_fd_sc_hd__dfbbn_1_3/Q_N FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0189f
C2285 FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_DFF17.Q 0.256f
C2286 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__nand3_1_2/Y 4.18e-19
C2287 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00246f
C2288 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_193_47# -0.0128f
C2289 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 8e-19
C2290 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_48/Y 9.5e-20
C2291 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# V_LOW -0.102f
C2292 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 6.18e-20
C2293 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 4.29e-20
C2294 sky130_fd_sc_hd__conb_1_20/LO V_LOW 0.149f
C2295 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.581f
C2296 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0039f
C2297 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__inv_16_41/Y 0.475f
C2298 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__conb_1_14/HI 6.65e-19
C2299 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 0.00262f
C2300 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0111f
C2301 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00112f
C2302 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 1.56e-20
C2303 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 2.92e-19
C2304 sky130_fd_sc_hd__inv_1_33/Y V_LOW 0.336f
C2305 sky130_fd_sc_hd__conb_1_21/HI V_LOW 0.193f
C2306 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# sky130_fd_sc_hd__conb_1_39/HI -1.79e-19
C2307 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 0.0011f
C2308 sky130_fd_sc_hd__conb_1_31/LO V_LOW 0.0787f
C2309 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0152f
C2310 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__inv_16_42/Y 0.00219f
C2311 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.0303f
C2312 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__conb_1_33/HI 3.29e-20
C2313 RISING_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0303f
C2314 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__conb_1_8/LO 0.0122f
C2315 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__inv_1_27/Y 0.00742f
C2316 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# Reset 0.00124f
C2317 sky130_fd_sc_hd__inv_1_34/Y V_LOW 0.19f
C2318 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI 7.57e-19
C2319 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# 0.00163f
C2320 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_24/A 0.256f
C2321 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__conb_1_31/HI 3e-19
C2322 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00385f
C2323 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 4.15e-20
C2324 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_24/LO 6.18e-19
C2325 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 5.1e-21
C2326 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 2.39e-20
C2327 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 0.00137f
C2328 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 5.41e-22
C2329 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00117f
C2330 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 8.52e-19
C2331 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/Q_N -9.56e-20
C2332 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_66/A 4.01e-19
C2333 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__conb_1_2/HI 0.00211f
C2334 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00106f
C2335 sky130_fd_sc_hd__inv_16_6/A FULL_COUNTER.COUNT_SUB_DFF0.Q 1.25f
C2336 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_16_42/Y 0.153f
C2337 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# sky130_fd_sc_hd__inv_1_59/Y 3.94e-21
C2338 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__conb_1_30/HI 3.22e-21
C2339 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.26e-19
C2340 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# -0.00774f
C2341 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# -0.00239f
C2342 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# -0.00901f
C2343 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1_13/LO 0.0116f
C2344 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 2.27e-20
C2345 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.00397f
C2346 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.15e-20
C2347 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00195f
C2348 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__conb_1_12/LO 7.49e-19
C2349 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_15/HI 2.67e-20
C2350 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00285f
C2351 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_31/LO 0.00134f
C2352 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# -6.8e-19
C2353 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# 3.23e-21
C2354 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# 6.31e-21
C2355 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# RISING_COUNTER.COUNT_SUB_DFF12.Q 7.36e-19
C2356 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# 6.52e-20
C2357 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__inv_1_40/Y 0.0158f
C2358 sky130_fd_sc_hd__inv_1_11/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00182f
C2359 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.08e-19
C2360 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_69/Y 0.0219f
C2361 V_SENSE sky130_fd_sc_hd__inv_1_61/Y 0.00129f
C2362 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1_26/HI 0.00256f
C2363 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/Q_N 0.0246f
C2364 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__nand2_1_5/Y 0.0179f
C2365 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.3e-19
C2366 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_581_47# -2.6e-20
C2367 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1_44/HI 1.47e-20
C2368 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 0.0123f
C2369 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.71e-19
C2370 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 0.0293f
C2371 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_1_21/Y 9.55e-19
C2372 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 0.0101f
C2373 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 2.03e-21
C2374 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0322f
C2375 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0181f
C2376 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_16_4/Y 0.00156f
C2377 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 9.38e-20
C2378 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 7.96e-20
C2379 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.57e-19
C2380 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 9.21e-20
C2381 sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 0.00119f
C2382 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 2.7e-20
C2383 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_48/Y 1.66f
C2384 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 1.32e-20
C2385 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# -3.86e-20
C2386 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# -0.00341f
C2387 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# V_LOW 0.0045f
C2388 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# V_LOW -4.4e-19
C2389 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# V_LOW 4.8e-20
C2390 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/Q_N 5.85e-22
C2391 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# -3.79e-20
C2392 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# -4.66e-20
C2393 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.27e-20
C2394 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# V_LOW 0.0121f
C2395 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_0/HI 0.0312f
C2396 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.83e-20
C2397 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_21/LO 3.72e-20
C2398 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# sky130_fd_sc_hd__inv_1_60/Y 0.00369f
C2399 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 0.0348f
C2400 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00706f
C2401 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# V_LOW 0.00855f
C2402 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# V_LOW -2.68e-19
C2403 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 3.92e-19
C2404 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 5.49e-21
C2405 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.58e-19
C2406 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00148f
C2407 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_31/Y 1.46e-19
C2408 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_791_47# 2.12e-19
C2409 sky130_fd_sc_hd__inv_1_67/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 7.95e-21
C2410 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_557_413# 2.87e-19
C2411 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# sky130_fd_sc_hd__inv_1_29/Y 2.91e-19
C2412 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 2.2e-20
C2413 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.83e-19
C2414 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.372f
C2415 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__conb_1_39/HI -2.17e-19
C2416 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_791_47# 1.15e-20
C2417 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.57e-19
C2418 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.0417f
C2419 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# sky130_fd_sc_hd__inv_1_9/Y 4.16e-21
C2420 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_67/A 0.235f
C2421 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# V_LOW 0.0256f
C2422 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# CLOCK_GEN.SR_Op.Q 1.07e-19
C2423 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 2.52e-21
C2424 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 9.03e-21
C2425 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 2.84e-20
C2426 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.33e-20
C2427 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0213f
C2428 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_381_47# 5.02e-19
C2429 sky130_fd_sc_hd__dfbbn_1_50/Q_N RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00877f
C2430 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_47/A 0.0118f
C2431 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_47/Y 0.0271f
C2432 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_59/Y 0.00922f
C2433 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.00127f
C2434 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.55e-19
C2435 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 9.68e-20
C2436 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 1.69e-19
C2437 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_581_47# -2.6e-20
C2438 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# sky130_fd_sc_hd__inv_1_32/Y 2.48e-20
C2439 sky130_fd_sc_hd__inv_1_33/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0587f
C2440 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_45/HI 0.0275f
C2441 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# V_LOW 0.00313f
C2442 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__inv_1_28/Y 0.0169f
C2443 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 4.5e-20
C2444 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/Q_N -4.33e-20
C2445 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 4.14e-20
C2446 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 1.29e-19
C2447 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_193_47# 0.00161f
C2448 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 0.0247f
C2449 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0114f
C2450 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 9.28e-19
C2451 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00109f
C2452 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00479f
C2453 sky130_fd_sc_hd__dfbbn_1_3/Q_N FULL_COUNTER.COUNT_SUB_DFF5.Q 8.97e-19
C2454 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0261f
C2455 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 0.00444f
C2456 sky130_fd_sc_hd__inv_1_54/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q 2.52e-21
C2457 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 0.00171f
C2458 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# -3.06e-20
C2459 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# -6.43e-20
C2460 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0548f
C2461 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__conb_1_39/LO 1.95e-20
C2462 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0492f
C2463 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__inv_1_36/Y 0.00102f
C2464 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# V_LOW 1.38e-19
C2465 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00162f
C2466 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# -1.06e-19
C2467 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0282f
C2468 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# sky130_fd_sc_hd__inv_16_41/Y 3.19e-19
C2469 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# sky130_fd_sc_hd__inv_1_59/Y 5.21e-19
C2470 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__conb_1_47/HI 1.05e-19
C2471 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_64/A 0.323f
C2472 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 2.57e-20
C2473 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_16/HI -0.0154f
C2474 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# -0.224f
C2475 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# -0.00419f
C2476 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__conb_1_28/HI 0.00305f
C2477 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# Reset 8.26e-19
C2478 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__inv_1_44/A 0.00267f
C2479 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# V_LOW 2.94e-20
C2480 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__inv_1_7/Y 1.19e-19
C2481 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.46e-19
C2482 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# V_LOW 0.0128f
C2483 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__nor2_1_0/Y 0.00281f
C2484 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00159f
C2485 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0226f
C2486 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_4/HI 1.59e-20
C2487 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# -0.00431f
C2488 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_473_413# -0.00458f
C2489 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 4.42e-20
C2490 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 4.42e-20
C2491 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 4.17e-20
C2492 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00136f
C2493 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 0.00384f
C2494 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 8.67e-19
C2495 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 1.38e-20
C2496 RISING_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 0.027f
C2497 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_0/a_27_47# 0.00153f
C2498 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# sky130_fd_sc_hd__inv_1_43/Y 3.62e-19
C2499 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 9.57e-20
C2500 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_24/Y 0.0015f
C2501 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# sky130_fd_sc_hd__inv_16_40/Y 0.00502f
C2502 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__conb_1_41/HI 2.61e-19
C2503 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00632f
C2504 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# -0.0014f
C2505 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# -7.89e-19
C2506 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00271f
C2507 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 4.38e-19
C2508 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 6.43e-20
C2509 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0396f
C2510 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.0156f
C2511 sky130_fd_sc_hd__dfbbn_1_27/Q_N RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00514f
C2512 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__inv_16_40/Y 0.0473f
C2513 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF17.Q -2.9e-20
C2514 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# V_LOW 0.0151f
C2515 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 7.27e-19
C2516 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.00125f
C2517 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.27e-20
C2518 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00403f
C2519 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.42e-19
C2520 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.239f
C2521 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_791_47# 4.27e-20
C2522 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 1.37e-20
C2523 sky130_fd_sc_hd__inv_1_37/Y V_LOW 0.378f
C2524 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_2/Y 0.0354f
C2525 RISING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.88e-20
C2526 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00541f
C2527 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# V_LOW 3.45e-19
C2528 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_66/Y 0.102f
C2529 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.93e-19
C2530 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 7.63e-19
C2531 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# V_LOW 1.38e-19
C2532 sky130_fd_sc_hd__inv_1_65/A Reset 0.0116f
C2533 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__nand2_8_4/Y 4.08e-20
C2534 sky130_fd_sc_hd__inv_1_48/Y CLOCK_GEN.SR_Op.Q 0.112f
C2535 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# -0.0198f
C2536 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 4.04e-19
C2537 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__conb_1_37/HI 1.78e-21
C2538 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 6.43e-19
C2539 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.493f
C2540 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 0.0141f
C2541 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__conb_1_47/HI 0.0347f
C2542 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00181f
C2543 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 5.18e-19
C2544 sky130_fd_sc_hd__inv_16_9/Y V_LOW 0.283f
C2545 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.012f
C2546 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 0.00429f
C2547 sky130_fd_sc_hd__conb_1_36/HI Reset 0.0836f
C2548 sky130_fd_sc_hd__conb_1_22/HI FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00126f
C2549 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# -3.57e-19
C2550 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# -3.86e-20
C2551 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0601f
C2552 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00278f
C2553 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_26/Y 0.155f
C2554 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__inv_1_35/Y 0.00438f
C2555 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0111f
C2556 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_14/LO 0.00643f
C2557 sky130_fd_sc_hd__conb_1_48/LO V_LOW 0.0825f
C2558 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# V_LOW 0.00306f
C2559 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.02e-21
C2560 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__conb_1_6/HI 2.66e-19
C2561 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# -1.44e-20
C2562 sky130_fd_sc_hd__conb_1_46/HI sky130_fd_sc_hd__conb_1_47/HI 0.0563f
C2563 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__conb_1_8/HI 0.00364f
C2564 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# sky130_fd_sc_hd__inv_1_7/Y 2.32e-20
C2565 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 3.92e-21
C2566 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# V_LOW 1.79e-20
C2567 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_1_21/Y 0.109f
C2568 sky130_fd_sc_hd__inv_1_66/A CLOCK_GEN.SR_Op.Q 0.0518f
C2569 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.00927f
C2570 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_20/Y 0.14f
C2571 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__nand2_1_5/Y 1.05e-19
C2572 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00201f
C2573 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.00158f
C2574 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_58/Y 0.0239f
C2575 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__conb_1_34/HI 0.0012f
C2576 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0919f
C2577 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 3.78e-19
C2578 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/Q_N 3.21e-19
C2579 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_47/Y 0.0093f
C2580 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_193_47# 0.00318f
C2581 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_28/HI 3.12e-19
C2582 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# -7.17e-20
C2583 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# -1.76e-19
C2584 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00363f
C2585 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0174f
C2586 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_2_0/A 1.8e-20
C2587 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__conb_1_29/HI 0.00922f
C2588 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__conb_1_19/HI 7.99e-20
C2589 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__conb_1_30/HI 0.0047f
C2590 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00848f
C2591 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 0.00848f
C2592 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_32/Y 0.00354f
C2593 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00578f
C2594 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 9.11e-19
C2595 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__inv_16_41/Y 3.57e-20
C2596 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__conb_1_21/HI 0.00398f
C2597 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 4.41e-19
C2598 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# 0.0109f
C2599 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 3.26e-19
C2600 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.12e-19
C2601 V_SENSE sky130_fd_sc_hd__inv_16_42/Y 0.00933f
C2602 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 4.24e-19
C2603 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_31/Y 1.26e-20
C2604 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_791_47# 4.01e-20
C2605 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_4_0/A 0.00816f
C2606 V_SENSE sky130_fd_sc_hd__conb_1_49/LO 9.19e-19
C2607 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.19e-20
C2608 RISING_COUNTER.COUNT_SUB_DFF13.Q V_LOW 1.81f
C2609 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 1.44e-19
C2610 sky130_fd_sc_hd__dfbbn_1_0/Q_N V_LOW -0.00135f
C2611 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_64/A 1.47e-21
C2612 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.99e-21
C2613 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_1_2/A 6.53e-19
C2614 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_61/Y 7.53e-21
C2615 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_1_22/Y 8.7e-19
C2616 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__inv_1_62/Y 5.54e-19
C2617 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_48/Y 4.14e-20
C2618 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# V_LOW -0.00266f
C2619 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00485f
C2620 sky130_fd_sc_hd__dfbbn_1_24/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 0.00185f
C2621 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# sky130_fd_sc_hd__conb_1_47/HI 4.97e-19
C2622 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 4.19e-20
C2623 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/Q_N 0.0327f
C2624 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__conb_1_25/HI -2.66e-19
C2625 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.36e-19
C2626 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0.0112f
C2627 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# -2.57e-20
C2628 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_16_41/Y 0.0203f
C2629 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0237f
C2630 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_29/Y 0.0708f
C2631 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__conb_1_38/HI 0.0581f
C2632 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 1.55e-20
C2633 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_25/Y 4.43e-21
C2634 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# V_LOW 0.00213f
C2635 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_51/Y 1.86e-19
C2636 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# -2.52e-19
C2637 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -0.00122f
C2638 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# V_LOW -2.78e-35
C2639 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_26/Y 8.32e-20
C2640 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__inv_1_41/Y 3.75e-21
C2641 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# sky130_fd_sc_hd__conb_1_5/HI 5.66e-21
C2642 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_58/Y 0.00778f
C2643 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# sky130_fd_sc_hd__conb_1_8/HI 0.00165f
C2644 sky130_fd_sc_hd__inv_16_50/Y V_SENSE 0.105f
C2645 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# sky130_fd_sc_hd__conb_1_23/HI 4.16e-19
C2646 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__inv_1_13/Y 1.22e-20
C2647 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_3/LO 4.45e-20
C2648 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# -2.32e-19
C2649 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# -0.00146f
C2650 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00136f
C2651 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_66/A 6.76e-22
C2652 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__conb_1_35/HI 3.34e-20
C2653 sky130_fd_sc_hd__dfbbn_1_3/Q_N FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0041f
C2654 sky130_fd_sc_hd__inv_1_11/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0333f
C2655 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# V_LOW 0.0576f
C2656 sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0776f
C2657 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__conb_1_34/HI -1.63e-19
C2658 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00173f
C2659 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__conb_1_38/HI 7.41e-19
C2660 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00889f
C2661 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.0133f
C2662 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__inv_1_25/Y 0.00525f
C2663 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__conb_1_27/HI -0.00908f
C2664 sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0168f
C2665 FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 2.68e-20
C2666 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# -0.00335f
C2667 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_557_413# -0.0012f
C2668 sky130_fd_sc_hd__conb_1_8/LO RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00218f
C2669 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 9.79e-20
C2670 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.75e-20
C2671 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# -0.00242f
C2672 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# -4.5e-20
C2673 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0309f
C2674 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_44/A 3.56e-19
C2675 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_1_34/Y 0.0047f
C2676 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 9.63e-19
C2677 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 9.63e-19
C2678 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 9.59e-19
C2679 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.0119f
C2680 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 1.09e-19
C2681 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 0.00267f
C2682 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_29/Y 5.83e-20
C2683 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00199f
C2684 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 0.113f
C2685 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 1.74e-20
C2686 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# V_LOW 0.0182f
C2687 sky130_fd_sc_hd__nand2_1_5/a_113_47# V_LOW -1.78e-19
C2688 sky130_fd_sc_hd__inv_1_28/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 1.73e-20
C2689 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# 1.8e-19
C2690 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/Q_N 0.00115f
C2691 sky130_fd_sc_hd__conb_1_6/HI sky130_fd_sc_hd__inv_1_10/Y 0.0389f
C2692 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 8.49e-19
C2693 sky130_fd_sc_hd__nor2_1_0/a_109_297# CLOCK_GEN.SR_Op.Q 0.00197f
C2694 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__conb_1_2/HI 0.00871f
C2695 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.53e-20
C2696 sky130_fd_sc_hd__inv_1_19/A FULL_COUNTER.COUNT_SUB_DFF2.Q 3.35e-21
C2697 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0303f
C2698 sky130_fd_sc_hd__inv_1_43/Y V_LOW 0.0885f
C2699 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# sky130_fd_sc_hd__conb_1_24/HI 0.00135f
C2700 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__inv_1_38/Y 0.00417f
C2701 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 1.36e-20
C2702 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 1.36e-20
C2703 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 5.32e-20
C2704 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# Reset 0.00143f
C2705 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__nand2_8_4/Y 1.5e-19
C2706 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI 0.00104f
C2707 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_0/LO 0.0142f
C2708 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# 1.68e-21
C2709 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# V_LOW 0.00571f
C2710 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.00479f
C2711 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.00109f
C2712 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 9.28e-19
C2713 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__inv_1_3/Y 1.96e-19
C2714 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__inv_1_54/Y 0.00574f
C2715 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00831f
C2716 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_21/Y 0.0192f
C2717 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 6.35e-21
C2718 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.287f
C2719 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# sky130_fd_sc_hd__conb_1_25/HI -3.88e-20
C2720 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.0706f
C2721 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__conb_1_0/HI 2.5f
C2722 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0846f
C2723 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 0.00143f
C2724 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__conb_1_41/HI 9.82e-20
C2725 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 3.31e-19
C2726 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0367f
C2727 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF0.Q 5.15e-20
C2728 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.168f
C2729 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# sky130_fd_sc_hd__inv_16_40/Y 5.32e-20
C2730 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 0.00713f
C2731 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.00107f
C2732 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# -1.76e-19
C2733 sky130_fd_sc_hd__dfbbn_1_4/Q_N V_LOW -0.00245f
C2734 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 1.67e-21
C2735 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 4.34e-20
C2736 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 9.21e-20
C2737 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00558f
C2738 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 1.01e-20
C2739 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.00523f
C2740 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__inv_1_58/Y 7.78e-21
C2741 sky130_fd_sc_hd__inv_16_8/A sky130_fd_sc_hd__inv_16_8/Y 0.319f
C2742 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_891_329# -2.2e-20
C2743 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -4.1e-19
C2744 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# -5.16e-20
C2745 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -1.64e-19
C2746 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.66e-19
C2747 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_647_21# 0.00185f
C2748 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 5.48e-21
C2749 sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# V_LOW 2.94e-20
C2750 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 1.89e-19
C2751 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.01e-20
C2752 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.045f
C2753 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 1.39e-19
C2754 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 2.62e-19
C2755 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__conb_1_27/HI -9.73e-19
C2756 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__conb_1_38/HI 1.11e-20
C2757 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 7.97e-19
C2758 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_30/HI 1.22e-21
C2759 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# V_LOW 0.0174f
C2760 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# V_LOW 4.8e-20
C2761 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# -0.00813f
C2762 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.78e-20
C2763 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.83e-19
C2764 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__inv_1_7/Y 0.00549f
C2765 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0393f
C2766 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# -0.0109f
C2767 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# -0.00631f
C2768 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0882f
C2769 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_51/Y 9.67e-19
C2770 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__conb_1_11/HI 0.00737f
C2771 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0161f
C2772 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.335f
C2773 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF17.Q 2.98e-19
C2774 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__inv_1_26/Y 0.00696f
C2775 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_1_49/Y 0.00521f
C2776 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# V_LOW 0.00566f
C2777 sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16_51/Y 1.36e-19
C2778 sky130_fd_sc_hd__inv_16_51/A sky130_fd_sc_hd__inv_16_49/A 0.0066f
C2779 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 5.82e-23
C2780 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 8.08e-20
C2781 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00219f
C2782 FALLING_COUNTER.COUNT_SUB_DFF1.Q transmission_gate_9/GN 0.00504f
C2783 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00244f
C2784 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00293f
C2785 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__conb_1_37/HI 0.00529f
C2786 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.37e-19
C2787 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 1.42e-19
C2788 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__conb_1_51/HI 8.99e-19
C2789 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_17/HI 5.48e-19
C2790 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 0.00386f
C2791 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__conb_1_12/HI 1.02e-19
C2792 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_37/Y 0.0263f
C2793 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_4_0/A 0.324f
C2794 V_SENSE sky130_fd_sc_hd__inv_16_2/Y 0.0256f
C2795 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 6.9e-21
C2796 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0249f
C2797 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# Reset 3.93e-20
C2798 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF15.Q -3.24e-20
C2799 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# -3.8e-20
C2800 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# -2.6e-19
C2801 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# -5.54e-21
C2802 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# CLOCK_GEN.SR_Op.Q 2.06e-20
C2803 FULL_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0288f
C2804 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# 4.04e-19
C2805 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 9.54e-19
C2806 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.00108f
C2807 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 4.99e-19
C2808 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0154f
C2809 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.69e-20
C2810 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 3.48e-20
C2811 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 2.04e-22
C2812 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 0.00291f
C2813 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__inv_1_33/Y 0.00312f
C2814 sky130_fd_sc_hd__inv_1_56/A Reset 4.3e-19
C2815 FALLING_COUNTER.COUNT_SUB_DFF2.Q transmission_gate_9/GN 1.28e-20
C2816 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__conb_1_44/HI 0.00815f
C2817 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 8.59e-20
C2818 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 0.00272f
C2819 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0159f
C2820 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# -4.66e-20
C2821 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# -3.79e-20
C2822 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 1.86e-21
C2823 sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00147f
C2824 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# Reset 8.68e-19
C2825 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# -0.00607f
C2826 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_891_329# -2.2e-20
C2827 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.46e-19
C2828 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 4.99e-20
C2829 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.00906f
C2830 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0956f
C2831 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_557_413# -0.0012f
C2832 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# -0.00393f
C2833 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__inv_16_40/Y 4.71e-20
C2834 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.27e-19
C2835 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_64/Y 0.105f
C2836 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_53/Y 0.172f
C2837 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# -0.00385f
C2838 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# -1.42e-32
C2839 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_29/LO 2.69e-19
C2840 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 1.98e-21
C2841 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_18/A 0.00671f
C2842 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_9/Y 2.31e-20
C2843 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_581_47# 5.8e-19
C2844 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# 8.26e-21
C2845 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.71e-19
C2846 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 2.87e-19
C2847 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.0141f
C2848 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__conb_1_27/HI -2.17e-19
C2849 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__inv_1_12/Y 1.21e-19
C2850 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__inv_1_26/Y 0.083f
C2851 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# -6.23e-21
C2852 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# -0.00367f
C2853 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 3.87e-19
C2854 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# V_LOW -0.107f
C2855 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# V_LOW 5.15e-20
C2856 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__conb_1_46/HI -0.00115f
C2857 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# V_LOW 0.00572f
C2858 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0393f
C2859 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# -0.00107f
C2860 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__conb_1_5/HI 0.0018f
C2861 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 2.18e-19
C2862 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# 0.00138f
C2863 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_1_12/Y 2.92e-21
C2864 sky130_fd_sc_hd__conb_1_0/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0233f
C2865 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/Q_N -9.56e-20
C2866 sky130_fd_sc_hd__dfbbn_1_35/Q_N FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0154f
C2867 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.07e-19
C2868 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0013f
C2869 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 7.82e-19
C2870 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# V_LOW 0.012f
C2871 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0306f
C2872 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0021f
C2873 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__conb_1_45/HI 1.04e-20
C2874 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_2/a_113_47# 2.49e-19
C2875 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# sky130_fd_sc_hd__inv_1_26/Y 5.98e-19
C2876 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_1_49/Y 0.0458f
C2877 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_16_42/Y 0.477f
C2878 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 6.79e-20
C2879 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.26e-21
C2880 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 1.95e-20
C2881 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_891_329# 7.18e-20
C2882 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 8.22e-20
C2883 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.021f
C2884 sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# sky130_fd_sc_hd__conb_1_12/HI -2.65e-20
C2885 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00133f
C2886 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__inv_1_37/Y 0.00552f
C2887 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 3.94e-20
C2888 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_4_0/A 0.0379f
C2889 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.00253f
C2890 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI -4.14e-19
C2891 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 0.00209f
C2892 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_29/Y 6.28e-20
C2893 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# -9.32e-20
C2894 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# V_LOW 0.00103f
C2895 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.00114f
C2896 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0.0116f
C2897 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.00278f
C2898 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 4.03e-19
C2899 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0.0116f
C2900 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# -1.24e-20
C2901 V_SENSE sky130_fd_sc_hd__fill_4_189/VPB 0.0258f
C2902 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.16e-19
C2903 sky130_fd_sc_hd__nand2_8_2/a_27_47# CLOCK_GEN.SR_Op.Q 0.0241f
C2904 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# sky130_fd_sc_hd__conb_1_29/HI -2.65e-20
C2905 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.92e-21
C2906 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_45/Y 1.46e-20
C2907 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# sky130_fd_sc_hd__conb_1_26/HI 3.78e-20
C2908 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 0.00364f
C2909 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# sky130_fd_sc_hd__inv_1_50/Y 7.05e-19
C2910 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_67/A 1.31e-21
C2911 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.00149f
C2912 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# -0.0169f
C2913 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_557_413# -0.0012f
C2914 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__conb_1_44/HI 1.1e-19
C2915 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__conb_1_43/HI 4.38e-19
C2916 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_47/Y 0.17f
C2917 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0172f
C2918 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# -0.00539f
C2919 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_36/HI 1.26e-19
C2920 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 8.39e-20
C2921 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.56e-19
C2922 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.84e-19
C2923 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/Q_N 9.65e-21
C2924 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 1.97e-19
C2925 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0729f
C2926 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 3e-21
C2927 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.81e-19
C2928 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 8.11e-21
C2929 sky130_fd_sc_hd__conb_1_8/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 0.275f
C2930 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.64e-19
C2931 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__nand3_1_1/Y 1.27e-19
C2932 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.00975f
C2933 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# sky130_fd_sc_hd__inv_16_40/Y 5.67e-19
C2934 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00105f
C2935 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0577f
C2936 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__conb_1_16/LO 4.72e-20
C2937 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# -4.66e-20
C2938 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# -3.79e-20
C2939 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# -0.0426f
C2940 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_4/HI 5.3e-20
C2941 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.27e-20
C2942 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__conb_1_16/HI 3.29e-20
C2943 sky130_fd_sc_hd__dfbbn_1_33/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 0.00185f
C2944 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.0375f
C2945 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# V_LOW -9.94e-19
C2946 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# -5.54e-21
C2947 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 1.33e-19
C2948 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# sky130_fd_sc_hd__conb_1_46/HI -2.07e-19
C2949 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 5.01e-19
C2950 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_1_47/Y 1.16e-21
C2951 sky130_fd_sc_hd__nand3_1_0/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 9.87e-21
C2952 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0455f
C2953 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.0149f
C2954 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0644f
C2955 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_24/HI 1.59e-19
C2956 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_22/Y 9.58e-21
C2957 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 0.0308f
C2958 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__inv_1_29/Y 0.0377f
C2959 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# -0.0203f
C2960 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_557_413# -3.67e-20
C2961 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand2_8_9/A 0.332f
C2962 sky130_fd_sc_hd__nand2_1_2/A FULL_COUNTER.COUNT_SUB_DFF1.Q 1.46e-20
C2963 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 1.06e-19
C2964 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__conb_1_43/LO 8.84e-20
C2965 sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__inv_1_62/Y 2.37e-20
C2966 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__inv_1_49/Y 3e-22
C2967 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_56/Y 3.14e-19
C2968 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 0.0173f
C2969 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 0.029f
C2970 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 7.9e-19
C2971 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 1.62e-19
C2972 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 2.27e-19
C2973 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_63/Y 0.0225f
C2974 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 6.63e-19
C2975 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_1_19/Y 2.98e-19
C2976 sky130_fd_sc_hd__conb_1_51/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0348f
C2977 sky130_fd_sc_hd__conb_1_49/LO sky130_fd_sc_hd__inv_1_63/Y 0.0121f
C2978 sky130_fd_sc_hd__conb_1_5/HI V_LOW 0.241f
C2979 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00124f
C2980 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# sky130_fd_sc_hd__inv_1_44/A 0.00114f
C2981 sky130_fd_sc_hd__inv_16_50/Y CLOCK_GEN.SR_Op.Q 0.0279f
C2982 sky130_fd_sc_hd__inv_1_11/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 1.98e-20
C2983 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__conb_1_32/HI 1.63e-20
C2984 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 0.026f
C2985 sky130_fd_sc_hd__conb_1_46/LO sky130_fd_sc_hd__conb_1_46/HI 7.46e-19
C2986 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 4.84e-19
C2987 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__conb_1_8/HI 4.17e-20
C2988 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/Q_N -4.33e-20
C2989 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_581_47# -2.6e-20
C2990 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_1_59/Y 6.3e-19
C2991 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 7.69e-19
C2992 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0.00193f
C2993 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__conb_1_5/LO 0.012f
C2994 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 6.56e-19
C2995 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0.0359f
C2996 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# 0.00199f
C2997 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__conb_1_0/HI 0.342f
C2998 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0483f
C2999 sky130_fd_sc_hd__inv_16_29/A sky130_fd_sc_hd__inv_16_8/A 0.0027f
C3000 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__conb_1_21/HI 1.4e-19
C3001 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# V_LOW -0.0723f
C3002 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 2.54e-20
C3003 FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0384f
C3004 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# -5.42e-19
C3005 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 7e-19
C3006 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__inv_1_10/Y 6.05e-20
C3007 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# V_LOW 4.8e-20
C3008 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__conb_1_44/HI 1.09e-19
C3009 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__inv_1_45/Y 0.00696f
C3010 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.25e-19
C3011 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# V_LOW -0.00121f
C3012 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 8.14e-20
C3013 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00119f
C3014 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0329f
C3015 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00842f
C3016 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_9/A 0.108f
C3017 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.25e-19
C3018 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_64/Y 5.39e-20
C3019 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 9.58e-20
C3020 sky130_fd_sc_hd__inv_1_4/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0443f
C3021 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# V_LOW 0.0148f
C3022 sky130_fd_sc_hd__inv_1_55/Y Reset 1.67e-19
C3023 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF7.Q 0.466f
C3024 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# V_LOW 1.38e-19
C3025 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# 2.05e-21
C3026 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.99e-19
C3027 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00174f
C3028 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__conb_1_16/LO 3.81e-20
C3029 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_941_21# 0.0239f
C3030 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__inv_1_69/Y 1.07e-20
C3031 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00307f
C3032 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/Q_N 6.01e-21
C3033 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0131f
C3034 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_1_47/Y 1.94e-22
C3035 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_30/Y 0.0213f
C3036 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# V_LOW 3.56e-20
C3037 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_1_42/Y 6.69e-20
C3038 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.00928f
C3039 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_647_21# -0.00157f
C3040 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_35/LO 3.52e-20
C3041 sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_9/A 0.00176f
C3042 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__conb_1_28/HI -0.0119f
C3043 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.06e-20
C3044 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# -5.42e-19
C3045 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# sky130_fd_sc_hd__inv_1_29/Y 5.12e-19
C3046 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.25e-21
C3047 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 1.33e-19
C3048 sky130_fd_sc_hd__conb_1_47/HI V_LOW 0.119f
C3049 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__conb_1_45/HI 1.66e-19
C3050 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 0.0415f
C3051 sky130_fd_sc_hd__inv_1_67/A Reset 0.00498f
C3052 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__conb_1_19/LO 1.64e-20
C3053 RISING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.82e-21
C3054 sky130_fd_sc_hd__conb_1_44/LO V_LOW 0.0878f
C3055 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# sky130_fd_sc_hd__conb_1_5/HI 9.52e-19
C3056 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__inv_1_61/Y 4.92e-19
C3057 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 2.75e-20
C3058 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 4.16e-19
C3059 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# Reset 0.0438f
C3060 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 9.59e-22
C3061 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__conb_1_23/HI -6.12e-19
C3062 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_30/LO 0.00525f
C3063 sky130_fd_sc_hd__conb_1_33/LO V_LOW 0.0951f
C3064 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 0.0326f
C3065 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# -2.18e-19
C3066 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# -3.51e-19
C3067 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 2.39e-20
C3068 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_791_47# 8.44e-19
C3069 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# 9.13e-19
C3070 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__conb_1_3/HI 7.52e-21
C3071 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# sky130_fd_sc_hd__conb_1_8/HI 6.39e-20
C3072 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# -5.84e-19
C3073 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# -0.0103f
C3074 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_30/HI 0.0192f
C3075 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF15.Q 1.44e-20
C3076 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_19/A 0.449f
C3077 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__conb_1_19/HI 0.0702f
C3078 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 0.0012f
C3079 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_41/HI 0.00544f
C3080 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__inv_1_31/Y 0.00315f
C3081 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# sky130_fd_sc_hd__conb_1_21/HI 4.02e-21
C3082 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# V_LOW -2.68e-19
C3083 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__conb_1_45/HI 0.0205f
C3084 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 1.31e-20
C3085 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__conb_1_19/HI 8.96e-20
C3086 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__conb_1_16/LO 9.17e-19
C3087 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__conb_1_23/HI 2.74e-20
C3088 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__conb_1_11/HI 1.39e-19
C3089 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 6.13e-19
C3090 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 9.06e-20
C3091 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0354f
C3092 sky130_fd_sc_hd__dfbbn_1_48/Q_N FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00862f
C3093 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.00172f
C3094 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 6.17e-19
C3095 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.93e-21
C3096 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0091f
C3097 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_1_10/Y 0.0564f
C3098 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__conb_1_14/LO 1.18e-20
C3099 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# sky130_fd_sc_hd__conb_1_6/HI 0.00138f
C3100 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_381_47# -2.53e-20
C3101 sky130_fd_sc_hd__conb_1_36/HI FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0811f
C3102 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# 0.00241f
C3103 sky130_fd_sc_hd__conb_1_41/HI FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.93e-19
C3104 sky130_fd_sc_hd__inv_1_10/Y V_LOW 0.0353f
C3105 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_2_0/A 0.583f
C3106 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__conb_1_7/HI 0.00412f
C3107 FULL_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0242f
C3108 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__inv_1_29/Y 0.101f
C3109 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_2_0/A 0.001f
C3110 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.36e-19
C3111 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__conb_1_15/HI 1.26e-19
C3112 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/Q_N -4.24e-20
C3113 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 4.08e-20
C3114 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 4.84e-20
C3115 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.0228f
C3116 sky130_fd_sc_hd__conb_1_3/HI V_LOW 0.196f
C3117 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0167f
C3118 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 1.42e-20
C3119 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 1.8e-21
C3120 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 6.72e-21
C3121 sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.00183f
C3122 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_581_47# -2.6e-20
C3123 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0255f
C3124 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_16_4/Y 0.0072f
C3125 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.17e-19
C3126 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00119f
C3127 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 0.042f
C3128 sky130_fd_sc_hd__conb_1_36/HI FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0376f
C3129 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_23/LO 0.0141f
C3130 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 5.48e-21
C3131 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_1_61/Y 3.07e-19
C3132 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# V_LOW 0.0153f
C3133 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__conb_1_32/HI 2.73e-20
C3134 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_33/Y 0.177f
C3135 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_1_39/Y 5.19e-19
C3136 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_891_329# 3.29e-20
C3137 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0145f
C3138 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 9.49e-19
C3139 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 1.16e-21
C3140 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# V_LOW 3.56e-20
C3141 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# Reset 0.00828f
C3142 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00148f
C3143 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# CLOCK_GEN.SR_Op.Q 0.0133f
C3144 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# V_LOW 0.00989f
C3145 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# sky130_fd_sc_hd__conb_1_23/HI -0.00256f
C3146 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_24/A 5.42e-19
C3147 RISING_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 0.856f
C3148 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00266f
C3149 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_791_47# 0.0023f
C3150 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__inv_1_1/Y 1.39e-20
C3151 sky130_fd_sc_hd__inv_4_0/A V_LOW 0.24f
C3152 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0206f
C3153 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__inv_1_25/Y 0.00519f
C3154 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.586f
C3155 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.84e-19
C3156 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# -6.8e-19
C3157 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF14.Q 0.101f
C3158 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__inv_1_60/Y 0.00348f
C3159 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# -3.86e-20
C3160 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# -0.00443f
C3161 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__conb_1_30/HI 0.00534f
C3162 Reset sky130_fd_sc_hd__inv_1_45/Y 0.00398f
C3163 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_45/Y 0.00785f
C3164 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.00504f
C3165 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/Q_N 7.56e-19
C3166 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0417f
C3167 sky130_fd_sc_hd__dfbbn_1_50/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00319f
C3168 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# V_LOW 7.36e-19
C3169 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__inv_1_14/Y 0.0107f
C3170 sky130_fd_sc_hd__inv_1_4/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0118f
C3171 sky130_fd_sc_hd__conb_1_0/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0187f
C3172 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.0308f
C3173 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# sky130_fd_sc_hd__conb_1_45/HI 5.15e-20
C3174 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# 7.28e-19
C3175 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__conb_1_41/HI -0.00115f
C3176 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 3.39e-19
C3177 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__conb_1_4/HI 0.0179f
C3178 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__conb_1_11/HI 1.33e-19
C3179 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# 8.88e-20
C3180 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__inv_1_38/Y 0.0288f
C3181 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_64/A 0.00841f
C3182 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_27/HI 0.061f
C3183 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_19/HI 3.63e-20
C3184 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__conb_1_29/HI 8.83e-21
C3185 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# sky130_fd_sc_hd__inv_1_10/Y 3.94e-21
C3186 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.019f
C3187 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__conb_1_50/HI 0.00114f
C3188 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# -6.43e-20
C3189 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# -0.00988f
C3190 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 9.63e-20
C3191 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00101f
C3192 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# -1.44e-20
C3193 sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__inv_1_44/A 0.00155f
C3194 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__conb_1_47/HI 9.88e-19
C3195 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# sky130_fd_sc_hd__inv_1_28/Y 7.05e-19
C3196 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# sky130_fd_sc_hd__conb_1_7/HI 3.49e-21
C3197 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 5.91e-20
C3198 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__inv_1_69/Y 5.85e-22
C3199 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__inv_1_21/Y 6.61e-20
C3200 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_44/A 0.018f
C3201 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# Reset 1.26e-19
C3202 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_7/Y 0.0585f
C3203 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_22/Y 1.79e-20
C3204 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0278f
C3205 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# -2.53e-20
C3206 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 0.00738f
C3207 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 2.2e-20
C3208 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_2_0/A 0.0416f
C3209 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 3.6e-19
C3210 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -0.00183f
C3211 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -7.6e-19
C3212 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.26e-20
C3213 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_25/HI 4.96e-20
C3214 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 1.21e-20
C3215 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__inv_1_55/Y 0.0101f
C3216 sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00269f
C3217 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_52/A 0.181f
C3218 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_1_0/Y 0.183f
C3219 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 1.89e-19
C3220 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_67/A 7.19e-21
C3221 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 8.26e-21
C3222 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 1.99e-19
C3223 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1_11/HI 2.86e-20
C3224 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF12.Q 0.675f
C3225 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_10/HI 0.00106f
C3226 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.00323f
C3227 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 8.64e-20
C3228 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__conb_1_51/HI 0.516f
C3229 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 1.65e-20
C3230 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# V_LOW -5.09e-19
C3231 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_4/a_113_47# 5.85e-19
C3232 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__conb_1_39/HI 7.98e-21
C3233 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# CLOCK_GEN.SR_Op.Q 0.00149f
C3234 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# -0.00402f
C3235 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# -3.86e-20
C3236 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 3.12e-19
C3237 sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__conb_1_26/HI 1.07e-20
C3238 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.52e-19
C3239 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# V_LOW 0.00161f
C3240 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# V_LOW 6.3e-19
C3241 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_9/Y 9.29e-20
C3242 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/Q_N -4.78e-20
C3243 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_30/Y 1.33e-19
C3244 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0769f
C3245 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 3.17e-20
C3246 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__conb_1_3/HI 2.11e-19
C3247 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00632f
C3248 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_9/HI 7.85e-20
C3249 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__conb_1_30/HI 0.00215f
C3250 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# -9.41e-19
C3251 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.0321f
C3252 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 8.75e-19
C3253 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# V_LOW -0.00916f
C3254 sky130_fd_sc_hd__conb_1_19/HI V_LOW 0.026f
C3255 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__inv_1_8/Y 0.0108f
C3256 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__conb_1_41/HI -2.07e-19
C3257 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 0.00249f
C3258 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__inv_1_61/Y 0.0118f
C3259 sky130_fd_sc_hd__conb_1_28/HI V_LOW 0.241f
C3260 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_16_4/Y 0.156f
C3261 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__conb_1_4/HI 1.34e-19
C3262 sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__conb_1_11/HI 6.37e-19
C3263 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 6.35e-21
C3264 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__inv_1_38/Y 0.00388f
C3265 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 1.08e-20
C3266 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_47/Y 0.211f
C3267 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.45e-19
C3268 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# V_LOW 0.00215f
C3269 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 3.79e-20
C3270 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_1_67/A 0.0538f
C3271 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 4.84e-21
C3272 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.78e-20
C3273 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# sky130_fd_sc_hd__conb_1_47/HI 1.79e-19
C3274 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00444f
C3275 sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0878f
C3276 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_51/HI 2.52e-19
C3277 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0111f
C3278 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__conb_1_15/LO 3.14e-20
C3279 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__inv_1_33/Y 0.044f
C3280 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# -5.54e-21
C3281 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# -3.8e-20
C3282 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -2.18e-19
C3283 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 0.137f
C3284 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 9.49e-20
C3285 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__inv_1_44/A 0.0053f
C3286 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q -4.98e-20
C3287 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 5.38e-20
C3288 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF11.Q 3.27e-19
C3289 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# -0.00141f
C3290 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# V_LOW 9.67e-20
C3291 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 0.0398f
C3292 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__conb_1_6/HI 0.0208f
C3293 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 1.83e-19
C3294 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 2.85e-20
C3295 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.027f
C3296 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.85e-20
C3297 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00711f
C3298 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00256f
C3299 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.62e-19
C3300 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00418f
C3301 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_46/A 0.213f
C3302 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# sky130_fd_sc_hd__inv_1_55/Y 2.36e-19
C3303 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__inv_1_43/Y 6.31e-21
C3304 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 0.00194f
C3305 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__conb_1_8/HI -7.65e-19
C3306 sky130_fd_sc_hd__conb_1_25/HI V_LOW 0.129f
C3307 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 2.48e-19
C3308 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# -2.53e-20
C3309 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00715f
C3310 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# V_LOW 0.00328f
C3311 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00131f
C3312 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# -9.41e-19
C3313 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 5.28e-19
C3314 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# V_LOW -0.0266f
C3315 sky130_fd_sc_hd__inv_1_25/Y V_LOW 0.353f
C3316 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# V_LOW 2.94e-20
C3317 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.11e-20
C3318 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__inv_1_30/Y 1.35e-20
C3319 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF0.Q 4.58e-19
C3320 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00641f
C3321 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.41e-21
C3322 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.032f
C3323 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__conb_1_7/HI 4.47e-20
C3324 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.156f
C3325 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_46/A 2.34e-20
C3326 V_SENSE transmission_gate_9/GN 16.3f
C3327 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# V_LOW 0.0129f
C3328 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__conb_1_20/HI 1.01e-19
C3329 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 0.0183f
C3330 sky130_fd_sc_hd__inv_1_53/A V_LOW 0.0609f
C3331 sky130_fd_sc_hd__dfbbn_1_29/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 0.00101f
C3332 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# V_LOW -0.00266f
C3333 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__conb_1_37/HI 1.57e-21
C3334 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# V_LOW 1.79e-20
C3335 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__inv_1_35/Y 0.00196f
C3336 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_6/HI 0.00268f
C3337 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0583f
C3338 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_41/LO 1.47e-19
C3339 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.118f
C3340 RISING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0309f
C3341 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_66/A 0.0016f
C3342 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_24/Y 0.307f
C3343 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 4.53e-19
C3344 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__conb_1_38/HI 0.00205f
C3345 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# V_LOW -0.018f
C3346 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# V_LOW 2.94e-20
C3347 sky130_fd_sc_hd__conb_1_24/HI RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0499f
C3348 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.31e-20
C3349 sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0872f
C3350 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_4/HI 3.19e-19
C3351 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0261f
C3352 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0197f
C3353 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__conb_1_51/HI 2.43e-19
C3354 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# sky130_fd_sc_hd__conb_1_44/HI 6.2e-19
C3355 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# V_LOW -0.329f
C3356 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.169f
C3357 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# -9.32e-20
C3358 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_19/HI 3.79e-19
C3359 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# 0.00198f
C3360 sky130_fd_sc_hd__inv_1_4/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0146f
C3361 sky130_fd_sc_hd__inv_1_47/A V_LOW 1.37f
C3362 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0207f
C3363 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0432f
C3364 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00481f
C3365 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.00367f
C3366 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_24/A 0.0723f
C3367 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__inv_1_9/Y 0.0308f
C3368 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.02f
C3369 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_32/HI 0.0239f
C3370 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_24/LO 2.61e-19
C3371 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/Q_N -4.33e-20
C3372 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 8.48e-19
C3373 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 1.58e-19
C3374 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.96e-20
C3375 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.83e-19
C3376 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.0266f
C3377 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0345f
C3378 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__conb_1_38/HI 0.0116f
C3379 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# 0.00161f
C3380 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__conb_1_8/HI 1.11e-20
C3381 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_6/HI 6.58e-22
C3382 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 1.06e-20
C3383 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 3.01e-19
C3384 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 5.66e-20
C3385 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 1.18e-20
C3386 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1_16/LO 8.01e-21
C3387 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# -1.44e-20
C3388 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_557_413# -3.67e-20
C3389 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# -0.00311f
C3390 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_891_329# -2.46e-19
C3391 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 6.02e-21
C3392 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__conb_1_17/HI 1.34e-20
C3393 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# V_LOW -0.0132f
C3394 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_1_64/A 8.25e-21
C3395 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 1.98e-19
C3396 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 9.75e-19
C3397 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 2.52e-19
C3398 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 1.68e-19
C3399 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0214f
C3400 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# 8.79e-22
C3401 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# -0.00216f
C3402 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_381_47# -0.00367f
C3403 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00388f
C3404 sky130_fd_sc_hd__dfbbn_1_47/Q_N RISING_COUNTER.COUNT_SUB_DFF0.Q 0.024f
C3405 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# sky130_fd_sc_hd__conb_1_7/HI -2.65e-20
C3406 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_29/Y 0.0334f
C3407 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# V_LOW 1.79e-20
C3408 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_43/LO 0.0181f
C3409 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.27e-22
C3410 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_23/Y 3.3e-19
C3411 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# 0.0015f
C3412 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0298f
C3413 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0.0371f
C3414 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0472f
C3415 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_16_8/Y 1.91e-19
C3416 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00147f
C3417 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_28/Y 0.0986f
C3418 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0311f
C3419 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__conb_1_24/HI 0.00953f
C3420 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__conb_1_31/HI 0.00107f
C3421 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_20/LO 2.22e-20
C3422 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__nand2_8_9/A 7.34e-20
C3423 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.77e-21
C3424 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 3.81e-20
C3425 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.14e-19
C3426 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.83e-19
C3427 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_19/A 0.00846f
C3428 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__conb_1_50/HI 1.21e-19
C3429 sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_28/Y 3.48e-19
C3430 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_891_329# -2.46e-19
C3431 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# -0.0238f
C3432 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_557_413# -3.67e-20
C3433 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00241f
C3434 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 1.58e-21
C3435 sky130_fd_sc_hd__conb_1_46/LO V_LOW 0.081f
C3436 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# -0.00458f
C3437 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# -0.00431f
C3438 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 3.72e-20
C3439 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# V_LOW -0.0084f
C3440 sky130_fd_sc_hd__inv_1_25/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00373f
C3441 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 1.86e-20
C3442 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 3.11e-19
C3443 sky130_fd_sc_hd__dfbbn_1_26/Q_N FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.94e-19
C3444 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_45/Y 7.6e-20
C3445 sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__inv_1_48/Y 0.0662f
C3446 FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 4.86e-20
C3447 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 0.288f
C3448 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__conb_1_43/HI 7.79e-21
C3449 sky130_fd_sc_hd__dfbbn_1_37/Q_N RISING_COUNTER.COUNT_SUB_DFF1.Q 0.022f
C3450 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0353f
C3451 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 8.27e-20
C3452 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.62e-21
C3453 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__conb_1_51/HI 4.38e-20
C3454 sky130_fd_sc_hd__conb_1_24/LO V_LOW 0.0667f
C3455 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__conb_1_48/HI 0.00286f
C3456 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00237f
C3457 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/Q_N -4.78e-20
C3458 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 9.03e-19
C3459 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 8.95e-20
C3460 sky130_fd_sc_hd__inv_16_15/A sky130_fd_sc_hd__inv_16_32/Y 0.0281f
C3461 sky130_fd_sc_hd__conb_1_12/HI V_LOW 0.278f
C3462 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0125f
C3463 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# 5.75e-19
C3464 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0258f
C3465 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 0.0198f
C3466 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__nor2_1_0/Y 8.61e-21
C3467 sky130_fd_sc_hd__conb_1_35/LO V_LOW 0.15f
C3468 sky130_fd_sc_hd__inv_1_40/Y sky130_fd_sc_hd__conb_1_30/HI 2.77e-21
C3469 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__inv_1_28/Y 0.0269f
C3470 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0107f
C3471 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 0.0269f
C3472 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.0109f
C3473 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_16_40/Y 0.059f
C3474 sky130_fd_sc_hd__dfbbn_1_21/Q_N FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.5e-19
C3475 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -1.89e-19
C3476 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# -3.87e-19
C3477 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_557_413# 4.09e-19
C3478 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0196f
C3479 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.45e-20
C3480 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_1_0/Y 0.00361f
C3481 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# V_LOW -0.00121f
C3482 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0389f
C3483 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.29e-19
C3484 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# -0.00441f
C3485 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# 9.42e-19
C3486 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF15.Q 9.52e-19
C3487 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 1.8e-20
C3488 sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__conb_1_37/HI 8.59e-19
C3489 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 1.76e-19
C3490 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_791_47# 1.41e-20
C3491 sky130_fd_sc_hd__inv_1_38/Y V_LOW 0.239f
C3492 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 2.88e-19
C3493 sky130_fd_sc_hd__dfbbn_1_22/Q_N V_LOW -0.00509f
C3494 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__conb_1_35/HI 2.92e-19
C3495 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.65e-20
C3496 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__conb_1_40/HI -0.00692f
C3497 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 1.06e-19
C3498 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.44e-20
C3499 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 5.82e-19
C3500 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_46/HI 3.34e-20
C3501 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.355f
C3502 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.022f
C3503 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# V_LOW 0.0132f
C3504 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_64/A 0.308f
C3505 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_8/HI 2.7e-20
C3506 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# V_LOW 4.8e-20
C3507 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 2.01e-20
C3508 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_791_47# 4.71e-20
C3509 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0334f
C3510 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_891_329# -2.2e-20
C3511 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# -0.00751f
C3512 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.0116f
C3513 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.0116f
C3514 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 4.03e-19
C3515 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.00278f
C3516 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.00114f
C3517 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.13f
C3518 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_381_47# 2.8e-20
C3519 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 3.67e-20
C3520 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 1.05e-19
C3521 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 1.05e-19
C3522 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0379f
C3523 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 2.9e-19
C3524 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0186f
C3525 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 8.26e-20
C3526 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 5.32e-20
C3527 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 2.42e-20
C3528 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 4.76e-19
C3529 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 1.38e-20
C3530 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0.00334f
C3531 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_1_26/Y 0.116f
C3532 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.19e-19
C3533 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.0216f
C3534 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__conb_1_24/HI 4.06e-19
C3535 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_15/A 0.0147f
C3536 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_30/Y 0.143f
C3537 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_66/A 0.0642f
C3538 sky130_fd_sc_hd__conb_1_16/HI FULL_COUNTER.COUNT_SUB_DFF12.Q 4.45e-21
C3539 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 1.36e-19
C3540 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__nand3_1_2/Y 0.0185f
C3541 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0123f
C3542 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_27/HI 2.2e-19
C3543 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 0.00931f
C3544 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.5e-20
C3545 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__nand2_1_2/A 1.54e-19
C3546 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# -0.00499f
C3547 sky130_fd_sc_hd__dfbbn_1_19/a_557_413# V_LOW 3.56e-20
C3548 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# sky130_fd_sc_hd__conb_1_50/HI -0.00162f
C3549 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# sky130_fd_sc_hd__conb_1_9/HI 9.76e-19
C3550 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_1_64/A 1.94e-19
C3551 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00112f
C3552 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0214f
C3553 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 1.2e-20
C3554 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 4.55e-20
C3555 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.125f
C3556 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# FULL_COUNTER.COUNT_SUB_DFF6.Q 4.97e-20
C3557 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0464f
C3558 FALLING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 0.369f
C3559 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_33/Y 0.00229f
C3560 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__conb_1_13/LO 1.53e-19
C3561 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00415f
C3562 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 8.44e-22
C3563 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__inv_1_34/Y 1.75e-19
C3564 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.331f
C3565 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__conb_1_14/HI -0.0068f
C3566 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_66/A 5.89e-20
C3567 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_63/Y 0.0913f
C3568 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.67e-19
C3569 sky130_fd_sc_hd__conb_1_23/LO RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0108f
C3570 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 7.54e-21
C3571 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 4.25e-20
C3572 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 2.99e-20
C3573 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 8.62e-21
C3574 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 7.44e-19
C3575 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__conb_1_39/HI 7.93e-21
C3576 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_891_329# 0.00162f
C3577 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__inv_1_50/Y 3.11e-21
C3578 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 0.00113f
C3579 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_48/Y 1.98e-19
C3580 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# Reset 0.0405f
C3581 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_3/Y 0.00169f
C3582 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0.00466f
C3583 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_55/Y 0.0242f
C3584 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# -1.76e-19
C3585 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_1_33/Y 3.13e-23
C3586 FALLING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0477f
C3587 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0416f
C3588 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# -0.00141f
C3589 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_1/LO 0.0345f
C3590 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_2/HI 0.00661f
C3591 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# sky130_fd_sc_hd__inv_1_41/Y 2.87e-19
C3592 sky130_fd_sc_hd__conb_1_11/LO FULL_COUNTER.COUNT_SUB_DFF18.Q 6.05e-21
C3593 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__inv_1_10/Y 0.0227f
C3594 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 9.93e-21
C3595 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_1_59/Y 8.84e-20
C3596 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0123f
C3597 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 1.57e-19
C3598 sky130_fd_sc_hd__conb_1_24/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00133f
C3599 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__conb_1_35/HI -5.86e-20
C3600 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_7/Y 1.21e-21
C3601 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__conb_1_38/LO 9.26e-19
C3602 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# sky130_fd_sc_hd__conb_1_40/HI 2.47e-19
C3603 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.111f
C3604 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.26e-20
C3605 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 0.00358f
C3606 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__inv_1_46/A 4.97e-20
C3607 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# -2.32e-19
C3608 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# -0.00135f
C3609 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 2.84e-32
C3610 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -0.00117f
C3611 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# -4.5e-20
C3612 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_67/A 0.292f
C3613 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0675f
C3614 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_557_413# 4.16e-19
C3615 sky130_fd_sc_hd__nand3_1_1/Y Reset 5.57e-20
C3616 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__nand3_1_1/Y 0.003f
C3617 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# -3.46e-20
C3618 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00504f
C3619 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/Q_N -7.69e-20
C3620 sky130_fd_sc_hd__inv_1_55/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 4.87e-20
C3621 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# 1.38e-19
C3622 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00326f
C3623 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# -0.00458f
C3624 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# -0.00423f
C3625 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_33/HI 0.134f
C3626 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_2_0/A 5.59e-19
C3627 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__inv_1_3/Y 8.46e-19
C3628 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.54e-19
C3629 sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF17.Q 0.187f
C3630 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 0.00301f
C3631 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_791_47# 2.82e-19
C3632 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 7.66e-21
C3633 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__inv_1_26/Y 0.0339f
C3634 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.42e-21
C3635 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# V_LOW 4.8e-20
C3636 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_66/Y 0.00362f
C3637 sky130_fd_sc_hd__inv_16_32/Y sky130_fd_sc_hd__inv_16_8/Y 1.92e-20
C3638 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 9.76e-20
C3639 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# V_LOW 0.064f
C3640 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.00114f
C3641 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_581_47# -2.6e-20
C3642 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# -0.115f
C3643 V_SENSE sky130_fd_sc_hd__conb_1_41/HI 0.00188f
C3644 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_32/A 3.58e-20
C3645 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__conb_1_19/LO 2.46e-20
C3646 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.29e-20
C3647 sky130_fd_sc_hd__nand2_8_3/a_27_47# V_LOW -0.0117f
C3648 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 6.22e-22
C3649 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_27/HI 1.14e-20
C3650 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_1_64/A 6.02e-21
C3651 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_22/A 0.0654f
C3652 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# sky130_fd_sc_hd__conb_1_3/HI 9.76e-19
C3653 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_60/Y 0.0311f
C3654 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# sky130_fd_sc_hd__nand3_1_2/Y 1.31e-19
C3655 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00468f
C3656 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0459f
C3657 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_647_21# -1.24e-20
C3658 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_29/A 0.00159f
C3659 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF6.Q 4.44e-20
C3660 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0569f
C3661 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# V_LOW 0.00732f
C3662 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 2.86e-20
C3663 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.46e-20
C3664 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.0304f
C3665 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.03e-19
C3666 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# sky130_fd_sc_hd__inv_1_34/Y 5.8e-19
C3667 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__conb_1_20/HI 4.12e-20
C3668 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# sky130_fd_sc_hd__conb_1_14/HI -9.33e-19
C3669 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_647_21# 9.42e-19
C3670 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.19e-20
C3671 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0106f
C3672 sky130_fd_sc_hd__dfbbn_1_43/Q_N FALLING_COUNTER.COUNT_SUB_DFF6.Q 4.38e-19
C3673 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_26/A 0.172f
C3674 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# sky130_fd_sc_hd__conb_1_39/HI 1.66e-19
C3675 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0.00115f
C3676 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 2.51e-19
C3677 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 2.17e-20
C3678 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_8/LO 4.64e-19
C3679 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__inv_1_27/Y 0.00665f
C3680 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# Reset 6.35e-20
C3681 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__conb_1_23/HI 0.00114f
C3682 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# 5.07e-19
C3683 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 2.67e-20
C3684 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 2.73e-21
C3685 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_1_0/Y 6.01e-21
C3686 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.0476f
C3687 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_66/A 0.181f
C3688 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# sky130_fd_sc_hd__conb_1_2/HI 5.75e-19
C3689 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__inv_1_24/A 0.00108f
C3690 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__inv_1_59/Y 9.37e-21
C3691 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__conb_1_43/HI 5.18e-19
C3692 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__conb_1_30/HI 1.36e-20
C3693 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__conb_1_29/HI 7.93e-20
C3694 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/Q_N 5.94e-21
C3695 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -0.00415f
C3696 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# -0.00563f
C3697 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 1.56e-20
C3698 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00237f
C3699 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# -0.00458f
C3700 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# -0.00423f
C3701 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 3.69e-19
C3702 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__conb_1_35/HI -2.17e-19
C3703 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__conb_1_40/HI -3.26e-20
C3704 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.035f
C3705 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_16_41/Y 0.462f
C3706 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__conb_1_12/LO 1.85e-19
C3707 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# 0.00199f
C3708 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 6.16e-19
C3709 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# sky130_fd_sc_hd__inv_1_1/Y 2.56e-21
C3710 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# -1.64e-19
C3711 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00229f
C3712 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__inv_1_69/Y 0.014f
C3713 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.8e-19
C3714 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 6.8e-19
C3715 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00162f
C3716 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/Q_N 5.16e-19
C3717 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 5.16e-19
C3718 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 0.0304f
C3719 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00167f
C3720 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 5.55e-21
C3721 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 2.53e-20
C3722 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 6.18e-21
C3723 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 2.02e-22
C3724 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.89e-20
C3725 sky130_fd_sc_hd__nand3_1_0/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 9.35e-20
C3726 sky130_fd_sc_hd__conb_1_45/HI FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0706f
C3727 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.44e-20
C3728 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_15/LO 0.00832f
C3729 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 1.41e-21
C3730 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_1_18/A 3.67e-19
C3731 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# -7.93e-19
C3732 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# -0.0014f
C3733 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_32/Y 1.41e-20
C3734 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# V_LOW -0.11f
C3735 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# V_LOW 0.00124f
C3736 RISING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.106f
C3737 sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# V_LOW 2.94e-20
C3738 sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.00172f
C3739 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00992f
C3740 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# V_LOW 0.0117f
C3741 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 1.02e-19
C3742 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.91e-20
C3743 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# sky130_fd_sc_hd__inv_1_60/Y 3.21e-19
C3744 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_48/A 0.0686f
C3745 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.0159f
C3746 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.93e-20
C3747 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.0951f
C3748 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 4.39e-19
C3749 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_581_47# -2.6e-20
C3750 sky130_fd_sc_hd__inv_1_35/Y sky130_fd_sc_hd__conb_1_32/HI 1.99e-21
C3751 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# V_LOW 0.00573f
C3752 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# V_LOW -0.00163f
C3753 sky130_fd_sc_hd__nand2_8_8/A FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00138f
C3754 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# sky130_fd_sc_hd__inv_16_40/Y 6.76e-20
C3755 sky130_fd_sc_hd__dfbbn_1_1/a_581_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 9.58e-20
C3756 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__conb_1_32/LO 0.012f
C3757 FULL_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0335f
C3758 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__conb_1_14/HI 4.34e-19
C3759 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_44/A 0.00296f
C3760 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00516f
C3761 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_891_329# 8.4e-19
C3762 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__inv_1_40/Y 6.89e-19
C3763 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_1_58/Y 3.8e-20
C3764 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# 1.67e-21
C3765 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__inv_1_29/Y 1.04e-19
C3766 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.76e-19
C3767 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.449f
C3768 sky130_fd_sc_hd__inv_1_8/Y RISING_COUNTER.COUNT_SUB_DFF7.Q 9.15e-21
C3769 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.113f
C3770 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.91e-19
C3771 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# sky130_fd_sc_hd__inv_1_9/Y 2.62e-20
C3772 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.066f
C3773 sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0325f
C3774 sky130_fd_sc_hd__inv_2_0/A Reset 0.0263f
C3775 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00328f
C3776 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# V_LOW 0.0142f
C3777 sky130_fd_sc_hd__inv_16_40/Y V_LOW 5f
C3778 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# CLOCK_GEN.SR_Op.Q 2.76e-19
C3779 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.51e-21
C3780 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 8.66e-22
C3781 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 8.85e-21
C3782 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0211f
C3783 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_47/A 2.69e-19
C3784 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_20/Y 0.124f
C3785 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__inv_1_66/A 1.82e-20
C3786 V_SENSE sky130_fd_sc_hd__inv_16_29/Y 0.483f
C3787 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_46/A 6.86e-19
C3788 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 2.44e-20
C3789 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0.0017f
C3790 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 7.66e-21
C3791 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0.00231f
C3792 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__conb_1_30/HI 2.28e-21
C3793 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 0.00463f
C3794 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 3.84e-19
C3795 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# -9.41e-19
C3796 FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 0.026f
C3797 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__inv_1_32/Y 1.1e-20
C3798 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__conb_1_12/LO 4.61e-20
C3799 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# V_LOW 4.91e-19
C3800 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_48/Y 1.21f
C3801 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__inv_1_28/Y 0.00655f
C3802 RISING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.01e-21
C3803 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 1.81e-20
C3804 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 1.23e-20
C3805 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_31/Y 2.23e-20
C3806 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 4.57e-21
C3807 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 8.83e-19
C3808 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 5.03e-19
C3809 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 7.67e-19
C3810 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__conb_1_10/HI 0.0234f
C3811 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 7.25e-19
C3812 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_791_47# 0.00698f
C3813 sky130_fd_sc_hd__conb_1_0/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0281f
C3814 sky130_fd_sc_hd__fill_8_848/VPB V_LOW 0.797f
C3815 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__inv_1_27/Y 1e-19
C3816 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.016f
C3817 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 9.55e-21
C3818 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# -3.86e-20
C3819 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# -0.00442f
C3820 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 5.32e-21
C3821 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.88e-21
C3822 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__conb_1_39/LO 1.22e-19
C3823 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0379f
C3824 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0276f
C3825 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_8/Y 0.00159f
C3826 sky130_fd_sc_hd__dfbbn_1_44/a_557_413# V_LOW 3.56e-20
C3827 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__conb_1_31/HI 8.83e-21
C3828 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# -1.76e-19
C3829 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# -7.17e-20
C3830 sky130_fd_sc_hd__conb_1_15/HI V_LOW 0.158f
C3831 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# sky130_fd_sc_hd__inv_1_32/Y 1.01e-20
C3832 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# V_LOW -9.94e-19
C3833 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__conb_1_28/LO 0.00334f
C3834 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_44/A 1.24e-19
C3835 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0216f
C3836 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# sky130_fd_sc_hd__inv_1_59/Y 9.76e-19
C3837 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_48/Y 0.0942f
C3838 sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16_55/Y 6.93e-19
C3839 sky130_fd_sc_hd__inv_16_51/A sky130_fd_sc_hd__inv_16_51/Y 0.0772f
C3840 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# -6.29e-19
C3841 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_891_329# -2.46e-19
C3842 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_557_413# -3.67e-20
C3843 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_16/HI -0.00125f
C3844 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# -0.0079f
C3845 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# Reset 0.0013f
C3846 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# sky130_fd_sc_hd__inv_1_44/A 7.46e-19
C3847 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.26e-20
C3848 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# 0.00203f
C3849 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__inv_1_7/Y 0.00839f
C3850 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 9.39e-20
C3851 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# V_LOW 0.0318f
C3852 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# sky130_fd_sc_hd__nor2_1_0/Y 4.94e-19
C3853 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00919f
C3854 sky130_fd_sc_hd__dfbbn_1_24/Q_N RISING_COUNTER.COUNT_SUB_DFF15.Q 4.52e-22
C3855 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 0.0429f
C3856 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_473_413# -0.012f
C3857 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# -0.00932f
C3858 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 4.99e-19
C3859 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 9.54e-19
C3860 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00108f
C3861 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__inv_1_58/Y 6.41e-22
C3862 sky130_fd_sc_hd__conb_1_33/HI FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.47e-21
C3863 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_0/a_193_47# 7.63e-21
C3864 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_34/HI 7.19e-19
C3865 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00743f
C3866 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# Reset 1.84e-20
C3867 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0173f
C3868 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# sky130_fd_sc_hd__inv_1_43/Y 1.49e-20
C3869 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__conb_1_12/LO 4.77e-21
C3870 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_30/LO 9.04e-21
C3871 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_1_6/Y 5.98e-20
C3872 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__inv_1_55/Y 1.42e-19
C3873 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__conb_1_41/HI 7.69e-19
C3874 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_1_39/Y 7.26e-19
C3875 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_1_24/Y 1.79e-19
C3876 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00149f
C3877 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# -0.00263f
C3878 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 5.68e-32
C3879 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -0.00226f
C3880 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__conb_1_30/HI 0.00519f
C3881 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 8.08e-21
C3882 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00634f
C3883 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.21e-20
C3884 sky130_fd_sc_hd__inv_1_14/Y V_LOW 0.143f
C3885 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 9.89e-21
C3886 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0303f
C3887 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 1.47e-20
C3888 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.00145f
C3889 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# V_LOW 0.00688f
C3890 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_791_47# 6.9e-19
C3891 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00612f
C3892 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.28e-19
C3893 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 1.19e-20
C3894 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 9e-19
C3895 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_1_66/Y 8.35e-20
C3896 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.74e-20
C3897 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_51/Y 0.26f
C3898 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0032f
C3899 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 1.32e-20
C3900 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# V_LOW 5.31e-20
C3901 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# sky130_fd_sc_hd__inv_1_28/Y 9.31e-20
C3902 sky130_fd_sc_hd__inv_16_15/Y sky130_fd_sc_hd__inv_16_28/Y 0.00529f
C3903 sky130_fd_sc_hd__inv_8_0/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00401f
C3904 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.38e-19
C3905 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# 1.22e-20
C3906 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 9.39e-19
C3907 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 2.02e-20
C3908 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# V_LOW 3.56e-20
C3909 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# -8.61e-20
C3910 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 1.61e-20
C3911 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# V_LOW 0.0164f
C3912 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0475f
C3913 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 0.0399f
C3914 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__conb_1_47/HI 0.0117f
C3915 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.32e-20
C3916 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# 1.93e-19
C3917 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 8.66e-20
C3918 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00328f
C3919 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__inv_1_30/Y 0.00511f
C3920 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# -9.41e-19
C3921 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# -7.77e-19
C3922 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# -2.15e-19
C3923 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.025f
C3924 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0417f
C3925 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 3.78e-19
C3926 sky130_fd_sc_hd__conb_1_18/LO V_LOW 0.0962f
C3927 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__conb_1_6/LO 0.00413f
C3928 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# sky130_fd_sc_hd__inv_1_35/Y 0.00147f
C3929 sky130_fd_sc_hd__inv_1_61/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.087f
C3930 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nand2_1_2/A 3.52e-20
C3931 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# V_LOW -0.00389f
C3932 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF15.Q 1.72e-20
C3933 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0167f
C3934 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__conb_1_16/HI -0.0127f
C3935 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_581_47# -7.91e-19
C3936 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 0.0246f
C3937 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_64/Y 0.0936f
C3938 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1_44/A 0.852f
C3939 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_16_2/Y 0.025f
C3940 sky130_fd_sc_hd__conb_1_29/LO V_LOW 0.0423f
C3941 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_8/HI 0.0162f
C3942 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.0013f
C3943 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 5.22e-20
C3944 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# V_LOW 0.0182f
C3945 sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 7.3e-20
C3946 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.0127f
C3947 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 7.53e-20
C3948 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_47/Y 2.22e-20
C3949 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# -2.57e-20
C3950 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 2.11e-19
C3951 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 6.38e-19
C3952 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# 2.11e-19
C3953 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# 6.38e-19
C3954 sky130_fd_sc_hd__nand2_1_3/a_113_47# V_LOW -1.78e-19
C3955 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__conb_1_34/HI -0.00543f
C3956 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.596f
C3957 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 1.16e-19
C3958 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/Q_N 9.65e-21
C3959 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 8.89e-20
C3960 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_19/LO 3.58e-20
C3961 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 4.52e-20
C3962 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__inv_1_6/Y 3.55e-19
C3963 V_SENSE sky130_fd_sc_hd__inv_1_56/A 5.01e-19
C3964 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 8.48e-19
C3965 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# -9.32e-20
C3966 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_2_0/A 2.43e-21
C3967 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_29/LO 1.8e-20
C3968 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__conb_1_19/HI 3.15e-21
C3969 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 4.19e-20
C3970 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_19/Y 0.0143f
C3971 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.12f
C3972 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_21/Y 3.77e-19
C3973 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.017f
C3974 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00185f
C3975 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.2e-20
C3976 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__conb_1_21/HI -4.9e-20
C3977 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.24e-19
C3978 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_1_31/Y 1.03e-20
C3979 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__inv_1_2/Y 3.97e-21
C3980 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__conb_1_40/HI 1.56e-20
C3981 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 2.76e-19
C3982 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 7.69e-20
C3983 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 3.13e-21
C3984 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_1_62/Y 5.93e-20
C3985 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 2.34e-20
C3986 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_42/Y 0.081f
C3987 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_581_47# -7.91e-19
C3988 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_48/Y 8.08e-19
C3989 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/Q_N 5.44e-19
C3990 sky130_fd_sc_hd__inv_1_65/A CLOCK_GEN.SR_Op.Q 0.0164f
C3991 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# V_LOW -6.55e-19
C3992 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.13e-19
C3993 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00486f
C3994 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# sky130_fd_sc_hd__conb_1_47/HI 1.16e-19
C3995 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_16_41/Y 2.31e-20
C3996 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_16_40/Y 5.12e-19
C3997 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__conb_1_25/HI -1.56e-20
C3998 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# -1.66e-19
C3999 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 8.2e-21
C4000 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.292f
C4001 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0278f
C4002 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_7/A 0.00124f
C4003 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 1.38f
C4004 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 8.9e-20
C4005 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# V_LOW 0.00398f
C4006 sky130_fd_sc_hd__conb_1_46/HI sky130_fd_sc_hd__inv_1_62/Y 8.04e-19
C4007 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -5.54e-21
C4008 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__inv_1_58/Y 7.04e-20
C4009 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# sky130_fd_sc_hd__conb_1_23/HI 0.00119f
C4010 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__nand2_8_8/A 1.51e-19
C4011 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# -0.00222f
C4012 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# -5.54e-21
C4013 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00225f
C4014 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__inv_1_13/Y 0.00107f
C4015 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__conb_1_35/HI 4.7e-20
C4016 sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.00148f
C4017 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_10/LO 4.18e-20
C4018 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# V_LOW 0.0123f
C4019 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# 0.0126f
C4020 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 7e-20
C4021 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__conb_1_38/HI 0.0041f
C4022 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0139f
C4023 sky130_fd_sc_hd__fill_8_951/VPB V_LOW 0.797f
C4024 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__inv_1_25/Y 0.00707f
C4025 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__conb_1_27/HI 0.00225f
C4026 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 7.69e-19
C4027 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__conb_1_34/HI -9.55e-19
C4028 V_SENSE sky130_fd_sc_hd__inv_16_48/A 0.554f
C4029 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0251f
C4030 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 2.57e-19
C4031 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_9/Y 3.37e-20
C4032 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# V_LOW 0.0589f
C4033 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# -0.00486f
C4034 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_891_329# -0.00159f
C4035 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_19/Y 0.00107f
C4036 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.05e-19
C4037 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# -0.00375f
C4038 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0199f
C4039 Reset V_LOW 2f
C4040 sky130_fd_sc_hd__nand2_8_4/Y V_LOW 0.115f
C4041 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/Q_N -4.78e-20
C4042 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__inv_1_13/Y 1.13e-19
C4043 sky130_fd_sc_hd__dfbbn_1_51/Q_N FALLING_COUNTER.COUNT_SUB_DFF10.Q 9.37e-20
C4044 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# sky130_fd_sc_hd__conb_1_19/HI 3.08e-21
C4045 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_1_34/Y 2.65e-21
C4046 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 0.00244f
C4047 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_28/Y 0.00345f
C4048 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_16_41/Y 0.192f
C4049 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 0.00244f
C4050 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.00599f
C4051 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.00132f
C4052 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.00142f
C4053 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 0.00105f
C4054 sky130_fd_sc_hd__conb_1_17/HI sky130_fd_sc_hd__inv_1_27/Y 4.97e-20
C4055 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.0157f
C4056 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# V_LOW 0.0137f
C4057 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_18/A 0.00689f
C4058 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0.00344f
C4059 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_24/A 0.00876f
C4060 sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 1.95e-19
C4061 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_39/LO 1.81e-20
C4062 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# sky130_fd_sc_hd__conb_1_21/HI -9.78e-19
C4063 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.94e-19
C4064 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 5e-20
C4065 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0262f
C4066 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.15e-20
C4067 sky130_fd_sc_hd__conb_1_51/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.053f
C4068 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_46/A 0.0277f
C4069 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.92e-19
C4070 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__conb_1_24/HI 5.83e-19
C4071 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 1.07e-20
C4072 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 1.07e-20
C4073 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_37/Y 6.14e-21
C4074 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# Reset 0.00101f
C4075 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__conb_1_30/HI 7.11e-20
C4076 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# V_LOW 0.011f
C4077 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 5.03e-19
C4078 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 7.67e-19
C4079 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 8.83e-19
C4080 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_1_48/Y 1.6e-19
C4081 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 6.34e-19
C4082 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__inv_1_3/Y 0.00198f
C4083 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.00109f
C4084 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_8/Y 0.089f
C4085 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.86e-20
C4086 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00237f
C4087 V_SENSE sky130_fd_sc_hd__inv_16_44/A 0.676f
C4088 sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 5.07e-19
C4089 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_41/HI 1.98e-19
C4090 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.023f
C4091 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_46/A 0.00349f
C4092 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# -0.0874f
C4093 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.708f
C4094 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 5.48e-21
C4095 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# V_LOW 1.79e-20
C4096 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__conb_1_4/HI 9.76e-19
C4097 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__conb_1_37/HI -7.59e-19
C4098 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 3.67e-21
C4099 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 8e-21
C4100 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 3.39e-20
C4101 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00116f
C4102 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 0.00803f
C4103 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 6.94e-19
C4104 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 5.52e-19
C4105 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__inv_1_58/Y 2.09e-21
C4106 V_SENSE sky130_fd_sc_hd__inv_16_7/Y 0.0159f
C4107 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# -4.66e-20
C4108 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -9.32e-20
C4109 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 8.38e-20
C4110 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_473_413# 0.00769f
C4111 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 1.33e-19
C4112 V_SENSE sky130_fd_sc_hd__inv_16_45/A 1f
C4113 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 6.28e-20
C4114 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0639f
C4115 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__conb_1_38/HI 6.59e-19
C4116 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 1.99e-20
C4117 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0.00784f
C4118 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 0.00987f
C4119 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00239f
C4120 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__conb_1_34/HI -1.58e-19
C4121 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# sky130_fd_sc_hd__conb_1_27/HI -6.57e-19
C4122 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0153f
C4123 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00567f
C4124 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF14.Q 2.03e-19
C4125 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nand2_8_8/A 0.32f
C4126 sky130_fd_sc_hd__inv_1_25/Y sky130_fd_sc_hd__conb_1_19/HI 0.00111f
C4127 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# V_LOW 0.0146f
C4128 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# V_LOW 2.94e-20
C4129 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# -3.46e-20
C4130 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# -0.0106f
C4131 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_557_413# -0.0012f
C4132 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_27_47# 0.0106f
C4133 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_14/HI 7.26e-22
C4134 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# -1.44e-20
C4135 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.44e-19
C4136 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# sky130_fd_sc_hd__inv_1_7/Y 1.82e-19
C4137 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0011f
C4138 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nand2_1_5/Y 1.87e-19
C4139 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# -0.0103f
C4140 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# -5.72e-19
C4141 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.53e-19
C4142 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 2.67e-19
C4143 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/Q_N 2.67e-19
C4144 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__conb_1_11/HI 0.00171f
C4145 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.0202f
C4146 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00454f
C4147 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 5.85e-20
C4148 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# sky130_fd_sc_hd__inv_16_41/Y 3.57e-20
C4149 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_1_26/Y 2.92e-19
C4150 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# V_LOW -5.05e-20
C4151 sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__inv_1_40/Y 1.41e-19
C4152 sky130_fd_sc_hd__inv_16_40/Y V_HIGH 2.08f
C4153 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__conb_1_10/HI 1.36e-20
C4154 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 5.58e-20
C4155 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_24/A 0.0234f
C4156 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 5.24e-19
C4157 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_14/LO 1.29e-19
C4158 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 1.63e-19
C4159 V_SENSE sky130_fd_sc_hd__inv_1_55/Y 5.42e-19
C4160 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00188f
C4161 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00441f
C4162 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# sky130_fd_sc_hd__conb_1_51/HI 2.11e-19
C4163 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 1.5e-19
C4164 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 6.55e-19
C4165 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# sky130_fd_sc_hd__conb_1_12/HI 5.03e-19
C4166 sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_56/Y 8.85e-19
C4167 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_1_37/Y 0.0208f
C4168 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_381_47# 0.0169f
C4169 sky130_fd_sc_hd__conb_1_46/HI FALLING_COUNTER.COUNT_SUB_DFF2.Q 1.59e-21
C4170 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0251f
C4171 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.00484f
C4172 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8_1/a_27_47# 0.0518f
C4173 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_8_9/A 0.0189f
C4174 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# -6.22e-19
C4175 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# -6.23e-21
C4176 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_381_47# -4.37e-20
C4177 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# V_LOW 1.79e-20
C4178 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0715f
C4179 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# 1.61e-20
C4180 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__inv_1_3/Y 1.54e-19
C4181 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_24/HI 2.43e-20
C4182 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 0.00942f
C4183 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 4.02e-19
C4184 sky130_fd_sc_hd__conb_1_49/LO FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.02e-19
C4185 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_24/A 5.66e-19
C4186 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.75e-21
C4187 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_19/A 0.0373f
C4188 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_581_47# 6.42e-19
C4189 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_2/Y 0.142f
C4190 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/Q_N 1.31e-19
C4191 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__conb_1_41/HI 3.05e-19
C4192 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__conb_1_44/HI 1.98e-19
C4193 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00352f
C4194 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0036f
C4195 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 3.05e-20
C4196 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 1.18e-20
C4197 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 8.26e-21
C4198 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.26e-19
C4199 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# Reset 0.00124f
C4200 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# -4.66e-20
C4201 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# -3.79e-20
C4202 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_1_38/Y 1.41e-20
C4203 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_25/Y 6.63e-21
C4204 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 4.72e-20
C4205 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.0122f
C4206 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/Q_N -4.78e-20
C4207 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 4.1e-19
C4208 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 5.86e-19
C4209 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00501f
C4210 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# 3.35e-19
C4211 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# -0.00524f
C4212 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_891_329# -0.00159f
C4213 sky130_fd_sc_hd__inv_1_44/A V_LOW 0.484f
C4214 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.29e-19
C4215 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_29/LO 1.14e-19
C4216 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__inv_1_28/Y 9.74e-20
C4217 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/Q_N -4.24e-20
C4218 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.06e-20
C4219 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# 5.98e-19
C4220 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_8/HI 9.19e-20
C4221 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_24/A 1.11e-19
C4222 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_36/Y 0.0684f
C4223 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# -0.116f
C4224 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_19/A 9.44e-22
C4225 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__conb_1_38/HI 8.96e-21
C4226 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0.0123f
C4227 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# 2.53e-19
C4228 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__conb_1_16/HI 0.0132f
C4229 sky130_fd_sc_hd__dfbbn_1_1/Q_N RISING_COUNTER.COUNT_SUB_DFF1.Q 2.83e-19
C4230 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.0371f
C4231 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 4.56e-20
C4232 FALLING_COUNTER.COUNT_SUB_DFF8.Q V_LOW 2.09f
C4233 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# -2.53e-20
C4234 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# V_LOW -0.00947f
C4235 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 0.00275f
C4236 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__conb_1_46/HI -0.00907f
C4237 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# V_LOW 0.0115f
C4238 sky130_fd_sc_hd__conb_1_24/HI FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.22f
C4239 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0412f
C4240 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 1.82e-20
C4241 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# -3.48e-19
C4242 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_647_21# 1.82e-19
C4243 sky130_fd_sc_hd__conb_1_22/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.2f
C4244 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__inv_1_12/Y 0.016f
C4245 sky130_fd_sc_hd__conb_1_21/HI RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0184f
C4246 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 3.46e-19
C4247 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00106f
C4248 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# -6.8e-19
C4249 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 5.66e-19
C4250 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# V_LOW 0.00738f
C4251 sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# sky130_fd_sc_hd__conb_1_11/HI -1.17e-19
C4252 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0312f
C4253 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 0.0354f
C4254 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 8.92e-20
C4255 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__conb_1_45/HI 0.00211f
C4256 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# sky130_fd_sc_hd__inv_1_49/Y 0.00125f
C4257 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_32/HI 5.18e-21
C4258 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 3.93e-20
C4259 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 8.25e-21
C4260 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00803f
C4261 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0163f
C4262 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# 1.07e-19
C4263 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0243f
C4264 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.48e-20
C4265 sky130_fd_sc_hd__dfbbn_1_31/a_581_47# sky130_fd_sc_hd__inv_1_37/Y 6.07e-19
C4266 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00125f
C4267 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 6.53e-19
C4268 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# -9.9e-19
C4269 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI -6.52e-20
C4270 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 1.88e-20
C4271 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# V_LOW 0.0125f
C4272 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_2/HI 0.00343f
C4273 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 1e-19
C4274 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 9.14e-19
C4275 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 7.34e-19
C4276 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# -3.06e-20
C4277 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# -6.43e-20
C4278 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/Q_N 5.44e-19
C4279 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 2.06e-20
C4280 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 5.31e-21
C4281 sky130_fd_sc_hd__inv_1_43/Y Reset 0.27f
C4282 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__inv_16_40/Y 0.444f
C4283 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 0.0171f
C4284 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_46/A 0.00426f
C4285 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# sky130_fd_sc_hd__conb_1_50/HI 6.1e-21
C4286 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# sky130_fd_sc_hd__inv_1_50/Y 2.78e-19
C4287 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_891_329# -0.00159f
C4288 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# -0.00548f
C4289 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_47/Y 1.53e-22
C4290 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 6.25e-21
C4291 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# V_LOW 0.043f
C4292 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# sky130_fd_sc_hd__conb_1_44/HI -2.65e-20
C4293 sky130_fd_sc_hd__inv_1_56/A CLOCK_GEN.SR_Op.Q 0.614f
C4294 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 2.42e-20
C4295 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00247f
C4296 sky130_fd_sc_hd__inv_1_68/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00458f
C4297 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_53/Y 5.51e-21
C4298 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00132f
C4299 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# CLOCK_GEN.SR_Op.Q 1.44e-19
C4300 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 9.97e-20
C4301 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 5.65e-19
C4302 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 0.00165f
C4303 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/Q_N 3.85e-20
C4304 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_48/LO 5.24e-19
C4305 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 5.62e-20
C4306 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00353f
C4307 sky130_fd_sc_hd__inv_16_31/Y V_LOW 0.164f
C4308 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0497f
C4309 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 1.18e-19
C4310 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 6.48e-20
C4311 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# -0.00385f
C4312 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00243f
C4313 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_29/LO 1.29e-19
C4314 sky130_fd_sc_hd__conb_1_38/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00161f
C4315 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 3.99e-20
C4316 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.72e-19
C4317 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00841f
C4318 sky130_fd_sc_hd__conb_1_13/HI FULL_COUNTER.COUNT_SUB_DFF15.Q 2.97e-21
C4319 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.57f
C4320 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_3/Y 6.64e-21
C4321 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.21e-19
C4322 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# -8.61e-20
C4323 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 2.32e-19
C4324 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00487f
C4325 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 0.00191f
C4326 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# -1.44e-20
C4327 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# V_LOW -0.00149f
C4328 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_381_47# -3.04e-19
C4329 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# -6.23e-21
C4330 sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__inv_1_38/Y 0.124f
C4331 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 7.52e-19
C4332 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__conb_1_46/HI -9.71e-19
C4333 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__inv_1_47/Y 2.88e-22
C4334 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00154f
C4335 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# V_LOW 1.79e-20
C4336 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 1.67e-21
C4337 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_24/HI 1.93e-19
C4338 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__inv_1_22/Y 0.0209f
C4339 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__conb_1_28/HI 0.0157f
C4340 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__inv_1_29/Y 0.0301f
C4341 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__inv_1_32/Y 0.00126f
C4342 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -0.00161f
C4343 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_891_329# -2.2e-20
C4344 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.00972f
C4345 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__conb_1_46/HI 1.17e-21
C4346 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q -2.16e-20
C4347 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 4.99e-21
C4348 sky130_fd_sc_hd__inv_1_63/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.326f
C4349 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__conb_1_38/HI 1.42e-20
C4350 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_1_49/Y 0.00575f
C4351 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00396f
C4352 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.73e-19
C4353 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI 0.0178f
C4354 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_29/A 0.0114f
C4355 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_5/HI 0.017f
C4356 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__conb_1_7/HI 0.00305f
C4357 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.00449f
C4358 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 6.25e-19
C4359 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 8.79e-21
C4360 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 4.81e-21
C4361 sky130_fd_sc_hd__conb_1_18/HI V_LOW 0.0192f
C4362 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_16_41/Y 0.00259f
C4363 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 1.14e-20
C4364 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_2_0/A 5.67e-19
C4365 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_51/A 0.151f
C4366 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 0.0121f
C4367 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00525f
C4368 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# sky130_fd_sc_hd__inv_1_44/A 0.00329f
C4369 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0305f
C4370 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00629f
C4371 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# -2.07e-19
C4372 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.94e-21
C4373 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# sky130_fd_sc_hd__conb_1_32/HI 6.43e-20
C4374 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 1.69e-19
C4375 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.86e-19
C4376 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 0.0505f
C4377 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# V_LOW 1.79e-20
C4378 sky130_fd_sc_hd__inv_1_64/Y V_LOW 0.0644f
C4379 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# sky130_fd_sc_hd__conb_1_25/HI 1.06e-21
C4380 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 6.57e-20
C4381 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0.0375f
C4382 sky130_fd_sc_hd__inv_16_48/A CLOCK_GEN.SR_Op.Q 0.0315f
C4383 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__conb_1_0/HI 0.0171f
C4384 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_1_33/Y 1.63e-21
C4385 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 2.4e-21
C4386 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_47/Y 6.18e-19
C4387 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# V_LOW 0.0193f
C4388 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# -3.46e-20
C4389 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__inv_1_10/Y 7.2e-20
C4390 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# V_LOW 2.94e-20
C4391 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0025f
C4392 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.257f
C4393 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__inv_1_45/Y 5.61e-19
C4394 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00231f
C4395 sky130_fd_sc_hd__conb_1_49/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.27e-20
C4396 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_56/A 1.05e-21
C4397 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# 2.57e-20
C4398 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# V_LOW -0.00266f
C4399 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.35e-20
C4400 sky130_fd_sc_hd__dfbbn_1_16/Q_N FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0373f
C4401 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0575f
C4402 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0174f
C4403 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 8.44e-21
C4404 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 4.19e-21
C4405 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_1_64/Y 8.77e-23
C4406 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00734f
C4407 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 0.0122f
C4408 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# V_LOW 0.0118f
C4409 sky130_fd_sc_hd__conb_1_51/HI FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0839f
C4410 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# V_LOW 3.56e-20
C4411 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_27_47# 0.229f
C4412 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 6.08e-21
C4413 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_11/Y 1.99e-21
C4414 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# 0.00226f
C4415 sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__nand3_1_1/Y 7.94e-20
C4416 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 0.00781f
C4417 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.7e-21
C4418 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_581_47# -7.91e-19
C4419 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__inv_1_69/Y 0.00611f
C4420 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_14/HI 5.23e-19
C4421 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__conb_1_46/HI -2.17e-19
C4422 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 5.74e-20
C4423 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.012f
C4424 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# V_LOW 2.26e-20
C4425 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_1_42/Y 5.54e-19
C4426 RISING_COUNTER.COUNT_SUB_DFF10.Q V_LOW 1.92f
C4427 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_647_21# -6.43e-20
C4428 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# -0.00932f
C4429 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_10/Y 0.0457f
C4430 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_891_329# 0.0014f
C4431 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__conb_1_24/HI 5.05e-19
C4432 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_60/Y 0.0236f
C4433 sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__inv_1_44/A 4.77e-20
C4434 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.26e-21
C4435 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__inv_1_29/Y 0.0555f
C4436 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# -3.46e-20
C4437 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_1_47/A 2.15e-19
C4438 sky130_fd_sc_hd__conb_1_49/LO sky130_fd_sc_hd__inv_1_60/Y 0.00108f
C4439 sky130_fd_sc_hd__conb_1_45/HI RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00266f
C4440 sky130_fd_sc_hd__inv_16_44/A CLOCK_GEN.SR_Op.Q 0.13f
C4441 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# 0.0385f
C4442 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__conb_1_45/HI 2.14e-20
C4443 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_16_41/Y 0.535f
C4444 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__conb_1_19/LO 9.91e-20
C4445 Reset V_HIGH 8.47f
C4446 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_3/HI 0.95f
C4447 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__conb_1_32/HI 0.00602f
C4448 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__conb_1_5/HI -2.07e-19
C4449 RISING_COUNTER.COUNT_SUB_DFF2.Q V_LOW 1.03f
C4450 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__inv_1_46/A 5.95e-19
C4451 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 2.69e-19
C4452 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 3.16e-19
C4453 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.43e-21
C4454 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_19/HI 0.00535f
C4455 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 6.98e-20
C4456 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# Reset 0.03f
C4457 sky130_fd_sc_hd__dfbbn_1_9/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00124f
C4458 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__conb_1_23/HI 0.0243f
C4459 FALLING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0199f
C4460 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_30/LO 0.00107f
C4461 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 0.00943f
C4462 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# -0.00117f
C4463 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# -9.88e-20
C4464 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# -0.00832f
C4465 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__conb_1_32/HI 1.38e-20
C4466 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_581_47# 2.34e-19
C4467 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# 0.00142f
C4468 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 3.84e-20
C4469 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# -2.52e-19
C4470 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# -0.00126f
C4471 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0134f
C4472 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_47/Y 0.0127f
C4473 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 9.17e-19
C4474 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF15.Q 1.04e-20
C4475 sky130_fd_sc_hd__inv_16_45/A CLOCK_GEN.SR_Op.Q 0.302f
C4476 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__conb_1_27/HI 1.89e-19
C4477 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_9/Y 2.85e-19
C4478 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_16_19/Y 4.6e-22
C4479 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__conb_1_0/HI 0.00241f
C4480 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_30/Y 1.15e-19
C4481 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_16_4/Y 2.05e-20
C4482 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.92e-21
C4483 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__inv_1_31/Y 3.44e-20
C4484 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/Q_N 1.47e-19
C4485 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# V_LOW 0.0127f
C4486 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/Q_N -6.48e-19
C4487 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00794f
C4488 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_24/Y 0.134f
C4489 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.94e-19
C4490 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_23/HI 0.00194f
C4491 sky130_fd_sc_hd__conb_1_18/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 5.23e-19
C4492 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__conb_1_50/HI 0.0024f
C4493 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.00251f
C4494 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 7.65e-21
C4495 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0359f
C4496 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0146f
C4497 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.01e-20
C4498 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0183f
C4499 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.84e-19
C4500 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_1_10/Y 0.00235f
C4501 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__conb_1_14/LO 3.07e-21
C4502 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00221f
C4503 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_557_413# -3.67e-20
C4504 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# -5.33e-20
C4505 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_14/LO 0.00251f
C4506 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__conb_1_51/HI 3.32e-20
C4507 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_2_0/A 0.0299f
C4508 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__conb_1_7/HI 0.00277f
C4509 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00178f
C4510 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 2.67e-20
C4511 sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 4.75e-19
C4512 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.61e-20
C4513 sky130_fd_sc_hd__inv_1_62/Y V_LOW 0.0441f
C4514 sky130_fd_sc_hd__conb_1_9/LO V_LOW 0.0493f
C4515 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.41e-21
C4516 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__conb_1_2/HI 0.02f
C4517 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0234f
C4518 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/Q_N -6.48e-19
C4519 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 3.46e-19
C4520 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# 0.0417f
C4521 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__conb_1_45/HI 7.4e-20
C4522 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00162f
C4523 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8_8/A 0.00639f
C4524 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_23/LO 0.00206f
C4525 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__conb_1_32/HI 4.52e-22
C4526 sky130_fd_sc_hd__inv_1_67/A CLOCK_GEN.SR_Op.Q 2.14e-19
C4527 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 1.33e-19
C4528 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# V_LOW 0.00241f
C4529 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_50/HI 0.508f
C4530 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 2.42e-19
C4531 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_53/A 2.26e-19
C4532 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# 1.13e-19
C4533 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 1.29e-20
C4534 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 2.93e-19
C4535 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.3e-20
C4536 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 3.39e-21
C4537 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# V_LOW 2.26e-20
C4538 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# Reset 2.17e-19
C4539 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00148f
C4540 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00186f
C4541 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__inv_1_33/Y 7.05e-20
C4542 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# CLOCK_GEN.SR_Op.Q 0.0297f
C4543 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# V_LOW 0.0122f
C4544 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_17/HI 4.31e-19
C4545 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_581_47# 6.57e-19
C4546 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__inv_1_1/Y 1.07e-20
C4547 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0226f
C4548 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0297f
C4549 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# 4.25e-20
C4550 sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__conb_1_8/HI 3.36e-20
C4551 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# -1.76e-19
C4552 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# sky130_fd_sc_hd__inv_1_60/Y 8.26e-19
C4553 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# -3.65e-19
C4554 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# -3.07e-19
C4555 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__conb_1_30/HI 2.43e-19
C4556 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_27/LO 8.52e-21
C4557 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.00439f
C4558 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.65e-20
C4559 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# V_LOW -0.102f
C4560 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.329f
C4561 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.0307f
C4562 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__conb_1_41/HI -0.00907f
C4563 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# 3.86e-19
C4564 sky130_fd_sc_hd__nor2_1_0/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0102f
C4565 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__conb_1_23/HI 6.57e-19
C4566 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.58e-21
C4567 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__conb_1_4/HI 0.00301f
C4568 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 4.76e-20
C4569 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 9.22e-20
C4570 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__inv_1_38/Y 0.0138f
C4571 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00116f
C4572 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00169f
C4573 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_19/HI 3.17e-19
C4574 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__conb_1_38/HI 5.62e-21
C4575 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_47/A 5.89e-20
C4576 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_29/HI 6.67e-20
C4577 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__inv_1_10/Y 9.37e-21
C4578 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0246f
C4579 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# sky130_fd_sc_hd__conb_1_50/HI 2.27e-19
C4580 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 0.36f
C4581 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# -9.35e-20
C4582 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# -3.86e-20
C4583 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 0.00333f
C4584 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00353f
C4585 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__conb_1_45/LO 1.48e-19
C4586 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_66/A 0.262f
C4587 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_47/HI 0.0362f
C4588 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__inv_1_28/Y 9.58e-19
C4589 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.29e-19
C4590 sky130_fd_sc_hd__conb_1_41/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 6.77e-20
C4591 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__conb_1_7/HI 0.00448f
C4592 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 1.83e-19
C4593 sky130_fd_sc_hd__conb_1_2/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00434f
C4594 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__inv_1_21/Y 1.16e-19
C4595 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__inv_1_13/Y 1.01e-19
C4596 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# Reset 3.22e-20
C4597 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_44/A 0.00649f
C4598 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 9.4e-19
C4599 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# -0.0163f
C4600 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_557_413# -3.67e-20
C4601 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 8.04e-21
C4602 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_15/HI 3.25e-19
C4603 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 6.18e-20
C4604 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0652f
C4605 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# -0.00472f
C4606 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -6.23e-21
C4607 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -6.22e-19
C4608 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__conb_1_25/HI 2.67e-20
C4609 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/Q_N 0.0263f
C4610 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 6.98e-20
C4611 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 1.64e-20
C4612 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__inv_1_55/Y 0.00238f
C4613 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 0.00153f
C4614 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__nand3_1_2/Y 1.26e-19
C4615 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_67/A 6.61e-19
C4616 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__inv_1_43/Y 1.85e-21
C4617 sky130_fd_sc_hd__conb_1_6/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00157f
C4618 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 5.79e-20
C4619 sky130_fd_sc_hd__nand2_8_9/Y V_LOW 0.0598f
C4620 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# V_LOW -0.106f
C4621 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# -2.66e-19
C4622 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# CLOCK_GEN.SR_Op.Q 4.19e-19
C4623 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# -2.28e-19
C4624 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.87e-20
C4625 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# V_LOW -0.115f
C4626 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# V_LOW 0.0163f
C4627 FALLING_COUNTER.COUNT_SUB_DFF1.Q V_LOW 1.3f
C4628 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_1_30/Y 4.19e-21
C4629 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 6.18e-20
C4630 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0257f
C4631 sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.403f
C4632 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.28e-20
C4633 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_9/HI 9.31e-20
C4634 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# -7.17e-20
C4635 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# -1.66e-19
C4636 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.036f
C4637 sky130_fd_sc_hd__dfbbn_1_17/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 6.48e-20
C4638 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# V_LOW 0.0463f
C4639 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# V_LOW 0.012f
C4640 sky130_fd_sc_hd__inv_1_45/Y CLOCK_GEN.SR_Op.Q 0.0121f
C4641 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# V_LOW -2.68e-19
C4642 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__inv_1_39/Y 0.00917f
C4643 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00307f
C4644 sky130_fd_sc_hd__conb_1_1/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 1.62e-19
C4645 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# sky130_fd_sc_hd__inv_16_40/Y 5.83e-21
C4646 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__conb_1_41/HI -9.71e-19
C4647 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 2.86e-20
C4648 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# sky130_fd_sc_hd__inv_1_38/Y 1.26e-19
C4649 FALLING_COUNTER.COUNT_SUB_DFF2.Q V_LOW 1.26f
C4650 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_8_0/Y 4.67e-20
C4651 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# sky130_fd_sc_hd__conb_1_19/HI 7.95e-20
C4652 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00658f
C4653 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 5.08e-20
C4654 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# -2.57e-20
C4655 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# V_LOW 0.0133f
C4656 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__conb_1_24/HI 1.8e-20
C4657 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# 4.36e-20
C4658 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 2.02e-19
C4659 sky130_fd_sc_hd__inv_1_39/Y V_LOW 0.379f
C4660 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# sky130_fd_sc_hd__conb_1_47/HI 7e-19
C4661 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 6.67e-22
C4662 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 8.79e-22
C4663 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__conb_1_51/HI 0.0226f
C4664 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00812f
C4665 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__conb_1_44/HI 0.00536f
C4666 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__conb_1_15/LO 2.6e-19
C4667 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 9.43e-20
C4668 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -9.88e-20
C4669 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# -6.23e-21
C4670 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# -4.37e-20
C4671 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.0543f
C4672 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 2.19e-19
C4673 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# sky130_fd_sc_hd__inv_1_44/A 2.41e-19
C4674 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# V_LOW -0.00551f
C4675 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.117f
C4676 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_1_3/Y 0.066f
C4677 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__conb_1_6/HI 9.77e-20
C4678 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 9.49e-20
C4679 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 6.76e-22
C4680 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.68e-19
C4681 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 2.68e-19
C4682 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00174f
C4683 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.015f
C4684 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 4.26e-19
C4685 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__inv_1_55/Y 6.42e-20
C4686 sky130_fd_sc_hd__inv_16_29/Y sky130_fd_sc_hd__inv_16_8/A 2.75e-19
C4687 V_SENSE sky130_fd_sc_hd__conb_1_46/HI 0.00178f
C4688 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0.00146f
C4689 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__conb_1_8/HI -0.0075f
C4690 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__inv_1_1/Y 0.109f
C4691 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_557_413# -3.67e-20
C4692 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# -0.00702f
C4693 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_891_329# -1.42e-19
C4694 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1_17/HI 1.18e-20
C4695 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 1.86e-21
C4696 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# V_LOW 1.38e-19
C4697 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# V_LOW -9.94e-19
C4698 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__conb_1_34/HI 1.36e-20
C4699 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1_31/HI 1.83e-19
C4700 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_17/HI 1.85e-20
C4701 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# -7.17e-20
C4702 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# -1.65e-19
C4703 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# V_LOW -0.00666f
C4704 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__conb_1_29/LO 5.12e-20
C4705 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00129f
C4706 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# V_LOW -2.68e-19
C4707 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0232f
C4708 sky130_fd_sc_hd__nand3_1_2/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 4.27e-19
C4709 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00158f
C4710 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 4.68e-21
C4711 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.55e-19
C4712 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0628f
C4713 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_33/Y 0.219f
C4714 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# V_LOW 0.0194f
C4715 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__conb_1_20/HI 1.55e-20
C4716 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 0.00807f
C4717 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_20/LO 4.53e-19
C4718 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00506f
C4719 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__conb_1_37/HI 1.98e-21
C4720 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# V_LOW -6.55e-19
C4721 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# V_LOW -0.00457f
C4722 FALLING_COUNTER.COUNT_SUB_DFF9.Q V_LOW 1.17f
C4723 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.559f
C4724 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__conb_1_41/HI -2.17e-19
C4725 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16_47/Y 0.00257f
C4726 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# 0.00178f
C4727 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 0.025f
C4728 sky130_fd_sc_hd__inv_16_6/A transmission_gate_9/GN 0.0864f
C4729 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.135f
C4730 sky130_fd_sc_hd__conb_1_2/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0877f
C4731 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 3.17e-21
C4732 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# V_LOW -0.00165f
C4733 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__inv_1_24/Y 1.15e-21
C4734 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__conb_1_36/LO 0.00525f
C4735 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00511f
C4736 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00301f
C4737 sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.94e-19
C4738 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0138f
C4739 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_21/LO 5.86e-21
C4740 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__conb_1_51/HI 4.96e-20
C4741 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.22e-19
C4742 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# sky130_fd_sc_hd__conb_1_44/HI 3.53e-19
C4743 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0947f
C4744 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_48/HI 0.0181f
C4745 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_8_8/A 3.38e-19
C4746 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# V_LOW -0.00991f
C4747 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 0.0577f
C4748 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 0.696f
C4749 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00886f
C4750 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0396f
C4751 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 9.23e-19
C4752 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.00238f
C4753 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0183f
C4754 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.56e-22
C4755 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.1e-20
C4756 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00869f
C4757 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__inv_16_40/Y 0.368f
C4758 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 0.00339f
C4759 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0223f
C4760 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_31/Y 0.0124f
C4761 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__conb_1_26/HI 0.0283f
C4762 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_16_41/Y 1.88e-20
C4763 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_18/A 0.00236f
C4764 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__conb_1_8/HI -9.48e-19
C4765 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 7.59e-20
C4766 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 9.68e-21
C4767 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 3.73e-19
C4768 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 8.63e-21
C4769 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# -4.36e-19
C4770 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_891_329# -3.3e-20
C4771 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# -0.00106f
C4772 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 1.17e-20
C4773 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 2.19e-20
C4774 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_50/A 0.212f
C4775 sky130_fd_sc_hd__conb_1_48/LO FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0483f
C4776 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 7.06e-21
C4777 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0107f
C4778 RISING_COUNTER.COUNT_SUB_DFF2.Q V_HIGH 1.89f
C4779 sky130_fd_sc_hd__dfbbn_1_8/Q_N FULL_COUNTER.COUNT_SUB_DFF14.Q 3.05e-19
C4780 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# V_LOW -1.39e-35
C4781 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_52/A 0.0241f
C4782 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# V_LOW 0.0642f
C4783 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 4.54e-19
C4784 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 6.66e-19
C4785 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 8.4e-21
C4786 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 0.003f
C4787 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 9.05e-19
C4788 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_381_47# -0.00375f
C4789 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.79e-19
C4790 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# 6.21e-21
C4791 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 8.31e-20
C4792 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# V_LOW 8.93e-19
C4793 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 4.24e-20
C4794 sky130_fd_sc_hd__dfbbn_1_19/a_1159_47# sky130_fd_sc_hd__conb_1_20/HI -1.05e-20
C4795 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_11/HI 2.65e-20
C4796 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.97e-19
C4797 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 1.97e-19
C4798 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.166f
C4799 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0249f
C4800 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__conb_1_0/HI 1.48e-19
C4801 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_47/A 5.25e-21
C4802 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0296f
C4803 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_20/LO 1.47e-19
C4804 sky130_fd_sc_hd__conb_1_4/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 1.02f
C4805 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.11e-20
C4806 sky130_fd_sc_hd__nand3_1_1/a_109_47# V_LOW -2.94e-19
C4807 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__nor2_1_0/Y 0.009f
C4808 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.52e-20
C4809 sky130_fd_sc_hd__inv_1_0/Y V_LOW 0.504f
C4810 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.34e-19
C4811 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00864f
C4812 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1_15/HI 4.39e-20
C4813 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__conb_1_50/HI -4.39e-19
C4814 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.366f
C4815 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_891_329# -2.2e-20
C4816 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# -0.00751f
C4817 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 1.81e-20
C4818 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 5.67e-19
C4819 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# -0.012f
C4820 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# -0.0126f
C4821 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.55e-20
C4822 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# V_LOW -1.39e-35
C4823 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 0.00108f
C4824 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00139f
C4825 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 9.87e-19
C4826 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_43/Y 0.267f
C4827 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__inv_1_39/Y 8.99e-21
C4828 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/Q_N -4.24e-20
C4829 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF7.Q 6.17e-19
C4830 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.18e-19
C4831 sky130_fd_sc_hd__nand2_8_8/A FULL_COUNTER.COUNT_SUB_DFF1.Q 7e-19
C4832 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00177f
C4833 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__conb_1_10/HI 3.8e-19
C4834 sky130_fd_sc_hd__conb_1_43/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.109f
C4835 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0526f
C4836 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# sky130_fd_sc_hd__conb_1_48/HI 8.82e-19
C4837 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.74e-19
C4838 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_0/a_113_47# 1.4e-19
C4839 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 4.12e-20
C4840 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 9.54e-19
C4841 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF9.Q 0.146f
C4842 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0416f
C4843 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_791_47# -0.0127f
C4844 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 1.93e-20
C4845 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 9.52e-20
C4846 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 9.52e-20
C4847 sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF17.Q 4.38e-19
C4848 sky130_fd_sc_hd__dfbbn_1_6/Q_N FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00264f
C4849 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# -0.00105f
C4850 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1_34/LO 0.0185f
C4851 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.28e-20
C4852 sky130_fd_sc_hd__inv_1_43/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 9.26e-22
C4853 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -2.18e-19
C4854 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# -2.01e-20
C4855 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_891_329# 3.43e-19
C4856 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__inv_1_0/Y 0.00275f
C4857 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00322f
C4858 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 0.0199f
C4859 FULL_COUNTER.COUNT_SUB_DFF18.Q V_LOW 3.01f
C4860 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# V_LOW -0.00266f
C4861 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00116f
C4862 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# 0.00395f
C4863 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00171f
C4864 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_557_413# -3.67e-20
C4865 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# -0.0209f
C4866 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__conb_1_51/HI 6.79e-19
C4867 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 4.5e-19
C4868 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__inv_1_14/Y 4.39e-19
C4869 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__conb_1_8/HI 8.96e-21
C4870 sky130_fd_sc_hd__inv_16_51/A sky130_fd_sc_hd__inv_16_55/Y 8.71e-19
C4871 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00738f
C4872 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# -0.00592f
C4873 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 2.88e-20
C4874 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_26/Y 9.4e-19
C4875 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__conb_1_35/HI 0.0205f
C4876 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_64/A 0.00684f
C4877 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__conb_1_40/HI 5.64e-19
C4878 sky130_fd_sc_hd__conb_1_42/HI V_LOW 0.0418f
C4879 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 9.19e-22
C4880 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 1.85e-22
C4881 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 8.98e-22
C4882 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.57e-19
C4883 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.0213f
C4884 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 5.01e-22
C4885 sky130_fd_sc_hd__dfbbn_1_43/Q_N V_LOW -0.0104f
C4886 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_46/HI 4.7e-20
C4887 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0194f
C4888 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0075f
C4889 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# V_LOW 0.00723f
C4890 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# V_LOW 2.94e-20
C4891 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_381_47# -3.79e-20
C4892 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# -4.66e-20
C4893 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0149f
C4894 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# -0.00141f
C4895 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# 1.3e-20
C4896 FALLING_COUNTER.COUNT_SUB_DFF12.Q V_LOW 1.46f
C4897 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 7.34e-19
C4898 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 9.14e-19
C4899 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 1e-19
C4900 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 0.0125f
C4901 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00234f
C4902 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00231f
C4903 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00233f
C4904 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 1.7e-20
C4905 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 4.64e-19
C4906 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 0.0107f
C4907 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 2.69e-19
C4908 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 0.00182f
C4909 RISING_COUNTER.COUNT_SUB_DFF14.Q V_LOW 1.43f
C4910 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_1_26/Y 0.0304f
C4911 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 8.03e-19
C4912 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00697f
C4913 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00101f
C4914 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_2/Y 0.0659f
C4915 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__conb_1_24/HI 2e-19
C4916 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# V_LOW 0.0158f
C4917 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_30/Y 0.0621f
C4918 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 7.17e-20
C4919 sky130_fd_sc_hd__inv_1_53/A Reset 4.82e-22
C4920 sky130_fd_sc_hd__nand2_8_4/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.11e-19
C4921 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 1.17e-20
C4922 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# -0.00122f
C4923 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# -0.00312f
C4924 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# V_LOW 2.26e-20
C4925 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# -3.46e-20
C4926 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__inv_1_64/A 1.58e-20
C4927 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__conb_1_39/HI 0.0018f
C4928 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# -2.57e-20
C4929 sky130_fd_sc_hd__dfbbn_1_49/Q_N V_LOW -0.0104f
C4930 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00188f
C4931 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 2.02e-20
C4932 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 8.11e-19
C4933 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0455f
C4934 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.29e-21
C4935 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nor2_1_0/Y 0.00464f
C4936 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0045f
C4937 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF6.Q 3.49e-19
C4938 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.3e-19
C4939 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_1_33/Y 5.44e-19
C4940 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__conb_1_37/HI 0.00513f
C4941 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.1e-19
C4942 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__inv_1_34/Y 0.00591f
C4943 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0206f
C4944 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__conb_1_14/HI 0.0017f
C4945 sky130_fd_sc_hd__inv_16_24/Y sky130_fd_sc_hd__inv_16_29/A 4.96e-19
C4946 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 7.57e-20
C4947 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_9/HI 4.01e-21
C4948 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_1_63/Y 2.96e-19
C4949 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 6.32e-19
C4950 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 7.51e-20
C4951 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 7.86e-20
C4952 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 1.26e-19
C4953 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 2.68e-20
C4954 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1_50/Y 0.0324f
C4955 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# 8.62e-19
C4956 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00882f
C4957 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# sky130_fd_sc_hd__inv_1_50/Y 0.00116f
C4958 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_24/Y 0.0228f
C4959 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# Reset 0.0348f
C4960 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# -2.07e-19
C4961 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 0.00868f
C4962 sky130_fd_sc_hd__conb_1_2/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00294f
C4963 sky130_fd_sc_hd__dfbbn_1_29/Q_N FALLING_COUNTER.COUNT_SUB_DFF6.Q 5.34e-22
C4964 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__inv_1_33/Y 8.34e-19
C4965 sky130_fd_sc_hd__inv_1_47/A Reset 0.0361f
C4966 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 0.00113f
C4967 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.283f
C4968 sky130_fd_sc_hd__inv_1_31/Y V_LOW 0.359f
C4969 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/Q_N 0.00188f
C4970 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# -5.42e-19
C4971 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_24/A 1.46e-19
C4972 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 0.00485f
C4973 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__nand2_1_5/Y 1.78e-19
C4974 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q -1.95e-19
C4975 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__inv_1_59/Y 0.00176f
C4976 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_29/HI 3.59e-19
C4977 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_24/HI 4.92e-19
C4978 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__inv_1_26/Y 6.58e-19
C4979 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__conb_1_35/HI 5.15e-20
C4980 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# sky130_fd_sc_hd__conb_1_40/HI -4.88e-19
C4981 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00576f
C4982 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 0.0354f
C4983 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.0348f
C4984 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0345f
C4985 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1_45/HI 1.38e-21
C4986 sky130_fd_sc_hd__conb_1_4/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 6.74e-19
C4987 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__inv_1_46/A 0.0011f
C4988 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# -2.02e-19
C4989 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# -5.54e-21
C4990 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# -0.00375f
C4991 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# sky130_fd_sc_hd__inv_1_49/Y 5.46e-20
C4992 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00277f
C4993 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0267f
C4994 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_891_329# 0.00119f
C4995 sky130_fd_sc_hd__inv_8_0/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00173f
C4996 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_51/A 9.14e-19
C4997 sky130_fd_sc_hd__conb_1_21/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0413f
C4998 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00341f
C4999 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# -0.012f
C5000 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -0.0037f
C5001 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_2_0/A 2e-19
C5002 FALLING_COUNTER.COUNT_SUB_DFF1.Q V_HIGH 1.75f
C5003 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_33/Y 0.0261f
C5004 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__inv_1_3/Y 0.00167f
C5005 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.68e-19
C5006 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_47/Y 8.72e-20
C5007 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_65/A 0.018f
C5008 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_26/HI 0.0171f
C5009 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 0.00425f
C5010 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 4.17e-20
C5011 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__inv_1_26/Y 7.69e-20
C5012 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.36e-20
C5013 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nand3_1_2/Y 0.239f
C5014 sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# V_LOW 2.94e-20
C5015 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# V_LOW 0.0189f
C5016 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_33/LO 0.00577f
C5017 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_24/A 8.63e-21
C5018 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# -0.00399f
C5019 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0994f
C5020 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.1e-21
C5021 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_60/Y 0.0283f
C5022 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_8/A 0.00136f
C5023 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# sky130_fd_sc_hd__nand3_1_2/Y 1.33e-19
C5024 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0031f
C5025 FALLING_COUNTER.COUNT_SUB_DFF2.Q V_HIGH 1.73f
C5026 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_647_21# -6.43e-20
C5027 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# -3.06e-20
C5028 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 7.14e-20
C5029 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00342f
C5030 FALLING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 1.35f
C5031 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 2.26e-19
C5032 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__inv_16_41/Y 0.0176f
C5033 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00185f
C5034 sky130_fd_sc_hd__dfbbn_1_24/a_581_47# sky130_fd_sc_hd__inv_1_33/Y 8.01e-20
C5035 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# V_LOW 0.00504f
C5036 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.0312f
C5037 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0713f
C5038 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00101f
C5039 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 0.0353f
C5040 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__conb_1_51/HI 0.102f
C5041 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# sky130_fd_sc_hd__conb_1_14/HI -6.57e-19
C5042 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_41/HI 0.0251f
C5043 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.53e-20
C5044 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_473_413# 0.0111f
C5045 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF1.Q 1.26e-19
C5046 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 8.84e-20
C5047 sky130_fd_sc_hd__dfbbn_1_42/a_581_47# sky130_fd_sc_hd__inv_1_63/Y 1.69e-19
C5048 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.113f
C5049 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__inv_16_41/Y 0.454f
C5050 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 4.42e-21
C5051 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 7.13e-21
C5052 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 0.281f
C5053 sky130_fd_sc_hd__conb_1_1/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 5.12e-21
C5054 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_1_63/Y 6.52e-20
C5055 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# 0.00211f
C5056 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__inv_16_41/Y 4.72e-19
C5057 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 2.55e-19
C5058 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 0.0013f
C5059 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 1.35e-19
C5060 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 3.43e-20
C5061 RISING_COUNTER.COUNT_SUB_DFF8.Q V_LOW 2.94f
C5062 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.38e-19
C5063 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# sky130_fd_sc_hd__conb_1_33/HI 2.13e-21
C5064 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_16_41/Y 0.0228f
C5065 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__inv_1_27/Y 0.00393f
C5066 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# Reset 0.00507f
C5067 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# CLOCK_GEN.SR_Op.Q 2.08e-20
C5068 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/Q_N -4.78e-20
C5069 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0.00346f
C5070 FULL_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0257f
C5071 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_36/HI 1.19e-20
C5072 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_1_66/A 8.46e-20
C5073 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__conb_1_2/HI 5.45e-20
C5074 sky130_fd_sc_hd__conb_1_46/HI sky130_fd_sc_hd__inv_1_63/Y 6.8e-19
C5075 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_19/Y 0.00546f
C5076 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__inv_1_24/A 8.32e-19
C5077 sky130_fd_sc_hd__conb_1_35/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 5.66e-20
C5078 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/Q_N 7.84e-20
C5079 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -0.0037f
C5080 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# -0.012f
C5081 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -4.39e-19
C5082 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# -2.52e-19
C5083 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_3/HI 5.93e-21
C5084 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.00179f
C5085 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_32/Y 0.182f
C5086 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__conb_1_25/HI 0.0042f
C5087 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# 1.84e-20
C5088 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 7.69e-20
C5089 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_18/LO 8.84e-20
C5090 sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00337f
C5091 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# -9.32e-20
C5092 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__inv_1_1/Y 6.8e-21
C5093 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# -0.00107f
C5094 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 3.6e-19
C5095 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# sky130_fd_sc_hd__inv_1_40/Y 6.1e-21
C5096 sky130_fd_sc_hd__nand3_1_1/Y CLOCK_GEN.SR_Op.Q 0.00132f
C5097 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00147f
C5098 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__inv_1_69/Y 6.24e-20
C5099 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.55e-19
C5100 V_SENSE sky130_fd_sc_hd__inv_16_50/A 0.367f
C5101 sky130_fd_sc_hd__dfbbn_1_29/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.79e-19
C5102 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# -2.57e-20
C5103 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0.00612f
C5104 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 0.238f
C5105 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_40/a_381_47# 0.00221f
C5106 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 0.0197f
C5107 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 0.00158f
C5108 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 9.08e-19
C5109 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 5.22e-22
C5110 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.47e-20
C5111 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 3.25e-19
C5112 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_1_26/Y 0.025f
C5113 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/Q_N 5.53e-19
C5114 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_31/Y 0.0913f
C5115 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__conb_1_32/HI 1.42e-21
C5116 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 6.25e-21
C5117 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 9.64e-19
C5118 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# -0.00226f
C5119 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# -0.00263f
C5120 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 2.47e-20
C5121 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# sky130_fd_sc_hd__inv_16_41/Y 7.11e-19
C5122 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# V_LOW -0.106f
C5123 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# V_LOW -0.0206f
C5124 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.0103f
C5125 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_581_47# -7.91e-19
C5126 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# V_LOW 0.00524f
C5127 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_67/A 3.19e-21
C5128 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 2.48e-19
C5129 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__inv_1_60/Y 0.00378f
C5130 sky130_fd_sc_hd__conb_1_2/LO RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0143f
C5131 sky130_fd_sc_hd__dfbbn_1_20/Q_N RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0291f
C5132 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_44/A 0.0324f
C5133 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.0725f
C5134 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00113f
C5135 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0013f
C5136 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_67/Y 0.0133f
C5137 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# V_LOW 0.0158f
C5138 sky130_fd_sc_hd__dfbbn_1_8/Q_N FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0339f
C5139 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_44/A 0.214f
C5140 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_15/HI 4.49e-19
C5141 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 0.00116f
C5142 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# sky130_fd_sc_hd__inv_16_40/Y 1.28e-19
C5143 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__conb_1_32/LO 5.65e-19
C5144 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__conb_1_19/HI 9.38e-20
C5145 sky130_fd_sc_hd__conb_1_50/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0899f
C5146 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.2e-19
C5147 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.0407f
C5148 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# 0.00256f
C5149 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00109f
C5150 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/Q_N 1.11e-19
C5151 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 3.67e-21
C5152 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 8e-21
C5153 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0425f
C5154 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_29/Y 0.379f
C5155 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00236f
C5156 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__inv_1_10/Y 0.0862f
C5157 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.24f
C5158 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0549f
C5159 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__inv_1_9/Y 3.3e-20
C5160 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.76e-19
C5161 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.587f
C5162 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 1.37e-19
C5163 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# sky130_fd_sc_hd__inv_1_27/Y 1.07e-21
C5164 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16_49/A 0.00341f
C5165 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# V_LOW 0.00908f
C5166 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.66e-20
C5167 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 7.58e-21
C5168 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 8.34e-20
C5169 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 2.11e-21
C5170 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.67e-19
C5171 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.013f
C5172 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_891_329# 0.00115f
C5173 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_47/A 4.26e-20
C5174 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 7.1e-19
C5175 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 8.73e-20
C5176 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 4.4e-20
C5177 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__inv_1_59/Y 6.01e-21
C5178 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 8.72e-19
C5179 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 0.00176f
C5180 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# -2.57e-20
C5181 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# -7.17e-20
C5182 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# -1.76e-19
C5183 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nand2_1_2/A 0.00115f
C5184 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_6/Q_N 3.58e-20
C5185 sky130_fd_sc_hd__dfbbn_1_26/Q_N FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0247f
C5186 sky130_fd_sc_hd__nand2_8_8/A FULL_COUNTER.COUNT_SUB_DFF0.Q 3.96e-20
C5187 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_1_28/Y 0.00174f
C5188 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__inv_16_40/Y 2.34e-19
C5189 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# V_LOW 3.56e-20
C5190 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/Q_N -4.24e-20
C5191 RISING_COUNTER.COUNT_SUB_DFF11.Q V_LOW 2.91f
C5192 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 2.18e-20
C5193 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# 1.28e-19
C5194 sky130_fd_sc_hd__conb_1_23/LO FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0567f
C5195 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 0.0035f
C5196 sky130_fd_sc_hd__inv_1_32/Y V_LOW 0.166f
C5197 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_24/A 0.00104f
C5198 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.0123f
C5199 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 1.66e-19
C5200 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__inv_1_36/Y 5.87e-21
C5201 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__inv_1_27/Y 5.36e-20
C5202 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0177f
C5203 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 1.25e-21
C5204 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# -3.65e-19
C5205 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# -3.07e-19
C5206 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 2.84e-32
C5207 V_SENSE V_LOW 33.3f
C5208 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 0.00167f
C5209 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 3.19e-22
C5210 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 7.69e-21
C5211 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__conb_1_44/LO 8.84e-20
C5212 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 0.026f
C5213 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.031f
C5214 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# V_LOW 2.26e-20
C5215 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# 3.59e-19
C5216 FALLING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.525f
C5217 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# -9.32e-20
C5218 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# V_LOW -9.94e-19
C5219 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# V_LOW 0.00283f
C5220 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__conb_1_27/HI 2.33e-20
C5221 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 5.63e-19
C5222 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00341f
C5223 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00911f
C5224 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_23/A 0.0019f
C5225 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 1.32e-19
C5226 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__conb_1_16/HI -0.00191f
C5227 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# -0.00431f
C5228 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# -0.0144f
C5229 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_891_329# -2.2e-20
C5230 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# -4.1e-19
C5231 sky130_fd_sc_hd__conb_1_4/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00588f
C5232 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__inv_1_44/A 9.33e-19
C5233 sky130_fd_sc_hd__conb_1_28/HI RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0022f
C5234 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 0.0259f
C5235 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_16_19/Y 0.00244f
C5236 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_1_7/Y 1.16e-19
C5237 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.3e-19
C5238 sky130_fd_sc_hd__dfbbn_1_39/Q_N V_LOW -0.00509f
C5239 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# V_LOW 0.00564f
C5240 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__conb_1_15/HI 0.00695f
C5241 sky130_fd_sc_hd__nand2_8_3/a_27_47# Reset 0.00341f
C5242 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# sky130_fd_sc_hd__nor2_1_0/Y 2.84e-20
C5243 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 2.14e-19
C5244 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 8.95e-22
C5245 sky130_fd_sc_hd__inv_16_41/Y V_LOW 1.57f
C5246 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 3.21e-21
C5247 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_1_44/A 2.29e-19
C5248 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# -0.0115f
C5249 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# -2.28e-19
C5250 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 6.72e-20
C5251 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 6.72e-20
C5252 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 0.00942f
C5253 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.49e-19
C5254 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF0.Q 3.45e-19
C5255 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 4.2e-20
C5256 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# Reset 7.69e-21
C5257 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0603f
C5258 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__conb_1_30/LO 9.25e-19
C5259 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__conb_1_41/HI 6.86e-21
C5260 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.3e-19
C5261 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 5.35e-20
C5262 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -0.00125f
C5263 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# -0.00472f
C5264 sky130_fd_sc_hd__inv_2_0/A CLOCK_GEN.SR_Op.Q 1.07e-19
C5265 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__conb_1_30/HI 5.85e-19
C5266 sky130_fd_sc_hd__nand2_8_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0526f
C5267 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.2e-19
C5268 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__inv_1_8/Y 0.013f
C5269 V_SENSE sky130_fd_sc_hd__inv_16_9/Y 0.046f
C5270 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.06e-20
C5271 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00637f
C5272 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_28/LO 0.0122f
C5273 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 4.15e-19
C5274 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# V_LOW 0.0163f
C5275 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.42e-20
C5276 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00289f
C5277 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__inv_16_41/Y 0.157f
C5278 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0021f
C5279 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 6.46e-20
C5280 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 9.58e-19
C5281 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00115f
C5282 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00136f
C5283 sky130_fd_sc_hd__conb_1_6/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 9.97e-20
C5284 sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0677f
C5285 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 8.06e-20
C5286 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_66/A 0.85f
C5287 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__nand2_1_5/Y 0.00104f
C5288 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 8.47e-21
C5289 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# V_LOW 2.26e-20
C5290 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_69/Y 5.68e-21
C5291 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__nand2_8_8/A 0.0108f
C5292 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_3/HI 0.184f
C5293 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# -0.0109f
C5294 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# -0.00631f
C5295 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 2.65e-20
C5296 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 5.05e-19
C5297 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# V_LOW -0.323f
C5298 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0462f
C5299 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.115f
C5300 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__conb_1_47/HI 0.0192f
C5301 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.41e-21
C5302 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00487f
C5303 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 8.81e-20
C5304 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# sky130_fd_sc_hd__inv_1_30/Y 8.39e-19
C5305 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_20/Y 0.0382f
C5306 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# -1.66e-19
C5307 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# -7.17e-20
C5308 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# -0.00183f
C5309 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00808f
C5310 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 0.00115f
C5311 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/Q_N -4.78e-20
C5312 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.46e-20
C5313 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# sky130_fd_sc_hd__inv_1_35/Y 1.45e-20
C5314 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 1.49e-19
C5315 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_16_42/Y 0.334f
C5316 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0015f
C5317 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 1.58e-19
C5318 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# V_LOW -9.15e-19
C5319 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00293f
C5320 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__conb_1_37/LO 8.81e-20
C5321 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# -0.00385f
C5322 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 0.0661f
C5323 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_5/HI 1.08e-20
C5324 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_3/HI 8.18e-22
C5325 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 1.21e-19
C5326 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_8/HI 0.011f
C5327 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.54e-20
C5328 FALLING_COUNTER.COUNT_SUB_DFF15.Q V_LOW 1.45f
C5329 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 1.34e-20
C5330 sky130_fd_sc_hd__inv_1_32/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.744f
C5331 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00778f
C5332 sky130_fd_sc_hd__inv_8_0/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 8.64e-20
C5333 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# -1.64e-19
C5334 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.032f
C5335 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 2.06e-20
C5336 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nor2_1_0/Y 3.85e-19
C5337 sky130_fd_sc_hd__conb_1_33/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.22e-21
C5338 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# Reset 9.3e-21
C5339 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_473_413# 5.17e-21
C5340 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__conb_1_28/HI 1.28e-20
C5341 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 7.83e-21
C5342 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_2_0/A 1.95e-20
C5343 sky130_fd_sc_hd__dfbbn_1_50/a_1159_47# sky130_fd_sc_hd__conb_1_30/HI 0.00183f
C5344 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_19/HI -0.0767f
C5345 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00404f
C5346 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00404f
C5347 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 5.63e-19
C5348 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.94e-21
C5349 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 3.25e-19
C5350 sky130_fd_sc_hd__dfbbn_1_24/a_581_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 3.32e-19
C5351 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.237f
C5352 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 0.00125f
C5353 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_66/Y 0.0037f
C5354 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# V_LOW 1.79e-20
C5355 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__conb_1_35/HI 0.0629f
C5356 sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 0.00137f
C5357 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_16_41/Y 0.0318f
C5358 sky130_fd_sc_hd__inv_16_40/Y Reset 0.447f
C5359 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_16_40/Y 3.57e-19
C5360 sky130_fd_sc_hd__nand2_8_0/a_27_47# V_LOW -0.00517f
C5361 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_24/HI 0.0155f
C5362 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.19e-20
C5363 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00463f
C5364 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 5.74e-20
C5365 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_4/HI 1.11e-20
C5366 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_9/HI 0.0747f
C5367 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_29/Y 2.57e-20
C5368 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 6.66e-20
C5369 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00612f
C5370 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_48/Y 5.04e-21
C5371 FULL_COUNTER.COUNT_SUB_DFF12.Q V_LOW 1.58f
C5372 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00379f
C5373 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_33/Y 1.1e-21
C5374 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.29e-20
C5375 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__conb_1_47/HI 0.00313f
C5376 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF15.Q 4.52e-22
C5377 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00122f
C5378 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__conb_1_25/HI -1.06e-20
C5379 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_44/A 1.13e-19
C5380 sky130_fd_sc_hd__conb_1_15/LO V_LOW 0.0352f
C5381 sky130_fd_sc_hd__conb_1_5/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00379f
C5382 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0957f
C5383 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.8e-20
C5384 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0117f
C5385 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# V_LOW 0.0147f
C5386 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -0.00117f
C5387 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_381_47# -0.00832f
C5388 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__inv_1_58/Y 0.00101f
C5389 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 1.14e-20
C5390 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_193_47# -0.0367f
C5391 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__conb_1_23/HI 0.00472f
C5392 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# -0.00216f
C5393 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# -4.5e-20
C5394 sky130_fd_sc_hd__dfbbn_1_7/Q_N V_LOW -0.00141f
C5395 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 9.59e-21
C5396 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__inv_1_13/Y 8.17e-22
C5397 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_35/HI 2.83e-20
C5398 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0222f
C5399 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# V_LOW 0.0153f
C5400 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 5.66e-19
C5401 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00199f
C5402 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/Q_N 5.66e-19
C5403 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_56/A 2.34e-19
C5404 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__conb_1_34/HI -6.57e-19
C5405 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__conb_1_38/HI 1.22e-20
C5406 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 9.4e-19
C5407 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_1_25/Y 0.00378f
C5408 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# sky130_fd_sc_hd__conb_1_27/HI 9.02e-19
C5409 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.00348f
C5410 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# sky130_fd_sc_hd__conb_1_20/HI 1.06e-21
C5411 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 0.00237f
C5412 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# V_LOW 0.0148f
C5413 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__inv_1_6/Y 1.87e-20
C5414 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# -0.00336f
C5415 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# -2.84e-32
C5416 sky130_fd_sc_hd__inv_16_50/A CLOCK_GEN.SR_Op.Q 0.0271f
C5417 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_33/Y 8.88e-19
C5418 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00219f
C5419 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q -3.24e-20
C5420 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__conb_1_27/HI 8.23e-22
C5421 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# -6.29e-19
C5422 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_557_413# -0.0012f
C5423 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_66/A 1.97e-20
C5424 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/Q_N -9.56e-20
C5425 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 0.00149f
C5426 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00149f
C5427 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_48/A 0.00192f
C5428 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 2.42e-19
C5429 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 1.08e-19
C5430 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.00109f
C5431 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# 8.63e-20
C5432 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 2.88e-19
C5433 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.00146f
C5434 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 8.18e-20
C5435 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0.0239f
C5436 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# V_LOW 0.00577f
C5437 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00281f
C5438 FALLING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 1.15e-19
C5439 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__conb_1_39/LO 2.37e-19
C5440 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_16_42/Y 0.113f
C5441 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0418f
C5442 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_10/Y 2.25e-19
C5443 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_16_41/Y 0.0207f
C5444 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# sky130_fd_sc_hd__inv_1_38/Y 5.46e-20
C5445 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_37/Y 2.14e-20
C5446 sky130_fd_sc_hd__inv_1_38/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00672f
C5447 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.22e-19
C5448 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# Reset 8.77e-19
C5449 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_1/Y 1.62e-20
C5450 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# V_LOW 0.0205f
C5451 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.0123f
C5452 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__inv_1_48/Y 4.71e-20
C5453 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__inv_1_3/Y 1.63e-19
C5454 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.58e-19
C5455 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.00996f
C5456 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.13e-19
C5457 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 0.00358f
C5458 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 7.23e-21
C5459 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__conb_1_47/HI 5.42e-19
C5460 sky130_fd_sc_hd__conb_1_48/HI V_LOW 0.124f
C5461 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# sky130_fd_sc_hd__conb_1_25/HI -2.92e-20
C5462 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_52/Y 0.0381f
C5463 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.0131f
C5464 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/Q_N -4.33e-20
C5465 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__conb_1_41/HI 2.08e-20
C5466 sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__conb_1_37/HI 2.43e-20
C5467 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00291f
C5468 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00438f
C5469 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 3.57e-19
C5470 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 5.21e-20
C5471 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_647_21# -8.61e-20
C5472 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.03f
C5473 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# Reset 0.0405f
C5474 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 1.33e-19
C5475 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.8e-20
C5476 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# -0.0501f
C5477 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 8.54e-19
C5478 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# V_LOW -0.00191f
C5479 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# sky130_fd_sc_hd__inv_1_25/Y 5.54e-20
C5480 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__conb_1_4/HI 0.0015f
C5481 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__conb_1_37/HI -7.62e-19
C5482 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 3.67e-20
C5483 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# 0.00416f
C5484 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 7.35e-19
C5485 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.00182f
C5486 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 5.79e-19
C5487 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.06e-21
C5488 sky130_fd_sc_hd__conb_1_43/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 3.22e-20
C5489 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_941_21# 3.82e-19
C5490 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.415f
C5491 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -3.04e-20
C5492 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.172f
C5493 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 3.1e-20
C5494 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 5.14e-19
C5495 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# sky130_fd_sc_hd__conb_1_38/HI 3.38e-19
C5496 sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.29e-19
C5497 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# sky130_fd_sc_hd__inv_1_25/Y 5.83e-21
C5498 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0016f
C5499 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 5.75e-19
C5500 sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__nand2_1_5/Y 0.336f
C5501 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_44/A 0.286f
C5502 sky130_fd_sc_hd__nand3_1_2/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.78e-20
C5503 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# V_LOW 0.00475f
C5504 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_18/HI 0.0108f
C5505 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_7/Y 1.16e-19
C5506 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_47/Y 0.0464f
C5507 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__inv_1_33/Y 9.52e-20
C5508 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_891_329# -0.00159f
C5509 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# -0.014f
C5510 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_193_47# 6.65e-19
C5511 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# -1.63e-19
C5512 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__nand2_1_5/Y 3.48e-20
C5513 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_2/Y 6.27e-20
C5514 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__conb_1_9/HI 1.23e-19
C5515 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# -0.00126f
C5516 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# -2.28e-19
C5517 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.23e-20
C5518 sky130_fd_sc_hd__inv_16_4/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.155f
C5519 CLOCK_GEN.SR_Op.Q V_LOW 1.49f
C5520 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_11/HI -0.0556f
C5521 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.23e-19
C5522 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 7.28e-21
C5523 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.0138f
C5524 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__inv_1_26/Y 1.5e-20
C5525 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# V_LOW -0.11f
C5526 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# sky130_fd_sc_hd__inv_1_45/Y 3.89e-19
C5527 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_1_50/Y 1.11e-19
C5528 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__conb_1_6/HI 2.05e-20
C5529 sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0576f
C5530 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.87e-19
C5531 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_64/Y 0.00221f
C5532 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 7.25e-19
C5533 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 2.14e-20
C5534 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_48/LO 0.00538f
C5535 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.19e-20
C5536 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.45e-20
C5537 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 0.00286f
C5538 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# sky130_fd_sc_hd__inv_1_10/Y 2.9e-20
C5539 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 1.25e-20
C5540 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_47/A 0.119f
C5541 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__conb_1_12/HI 0.00134f
C5542 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_557_413# 3.39e-19
C5543 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_1_37/Y 0.0151f
C5544 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.889f
C5545 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 2.58e-19
C5546 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__inv_1_37/Y 3.26e-20
C5547 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0229f
C5548 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 2.73e-20
C5549 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_381_47# -2.53e-20
C5550 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__conb_1_30/HI 1.86e-20
C5551 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_17/HI 4.04e-20
C5552 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# V_LOW 0.00591f
C5553 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 5.05e-19
C5554 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# 2.65e-20
C5555 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_1_48/Y 6.7e-20
C5556 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 2.38e-20
C5557 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 4.58e-19
C5558 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 7.44e-21
C5559 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0293f
C5560 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00134f
C5561 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0183f
C5562 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 0.00408f
C5563 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.49e-19
C5564 sky130_fd_sc_hd__inv_1_63/Y V_LOW 0.0647f
C5565 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 0.0245f
C5566 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# 7.13e-19
C5567 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 2e-21
C5568 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# sky130_fd_sc_hd__conb_1_41/HI 2.38e-19
C5569 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 9.26e-19
C5570 V_SENSE V_HIGH 9.97f
C5571 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 6.78e-19
C5572 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.144f
C5573 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__conb_1_16/HI 1.13e-22
C5574 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_581_47# -7.91e-19
C5575 sky130_fd_sc_hd__dfbbn_1_18/a_581_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.27e-19
C5576 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# Reset 7.85e-20
C5577 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 3.04e-19
C5578 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.45e-19
C5579 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__inv_1_38/Y 4.43e-21
C5580 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0201f
C5581 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 2.25e-19
C5582 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 2.4e-21
C5583 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 2.61e-19
C5584 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__conb_1_37/HI -0.0128f
C5585 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 5.63e-20
C5586 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 2.91e-19
C5587 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 1.95e-21
C5588 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# 4.57e-19
C5589 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# -0.00336f
C5590 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 4.23e-20
C5591 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 7.91e-21
C5592 sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_15/A 2.17e-20
C5593 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# 1.1e-19
C5594 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 0.0234f
C5595 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00354f
C5596 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.08e-20
C5597 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_29/LO 1.03e-20
C5598 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/Q_N -9.56e-20
C5599 FULL_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 1.73e-20
C5600 sky130_fd_sc_hd__conb_1_25/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.27e-21
C5601 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.21e-20
C5602 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00309f
C5603 sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 1.76e-19
C5604 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_36/Y 0.0289f
C5605 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 0.0012f
C5606 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# -0.00547f
C5607 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0176f
C5608 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00236f
C5609 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 9.18e-20
C5610 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.12f
C5611 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.0114f
C5612 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.83e-20
C5613 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_56/Y 1.54e-19
C5614 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 2.35e-20
C5615 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# -6.29e-19
C5616 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_557_413# -3.67e-20
C5617 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# V_LOW -0.00592f
C5618 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_557_413# 5.03e-19
C5619 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_52/A 5.67e-20
C5620 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__conb_1_46/HI 0.00105f
C5621 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0441f
C5622 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# V_LOW 0.0261f
C5623 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0164f
C5624 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# -0.00592f
C5625 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 3.55e-33
C5626 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__conb_1_5/HI 4.9e-20
C5627 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_791_47# 3.65e-19
C5628 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_473_413# 1.65e-20
C5629 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__conb_1_36/LO 9.51e-20
C5630 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.83e-19
C5631 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# -1.65e-19
C5632 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# V_LOW -0.108f
C5633 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_47/Y 0.00257f
C5634 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.166f
C5635 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00272f
C5636 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 3.2e-19
C5637 sky130_fd_sc_hd__dfbbn_1_18/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 0.00179f
C5638 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# V_LOW -9.94e-19
C5639 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.85e-20
C5640 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 1.14e-20
C5641 sky130_fd_sc_hd__dfbbn_1_4/Q_N FULL_COUNTER.COUNT_SUB_DFF12.Q 5.57e-20
C5642 sky130_fd_sc_hd__nand2_8_4/Y Reset 0.219f
C5643 sky130_fd_sc_hd__inv_1_30/Y V_LOW 0.108f
C5644 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# sky130_fd_sc_hd__inv_16_40/Y 1.3e-19
C5645 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.0431f
C5646 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0586f
C5647 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0036f
C5648 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# sky130_fd_sc_hd__inv_1_37/Y 7.27e-19
C5649 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 6.47e-20
C5650 sky130_fd_sc_hd__conb_1_46/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00667f
C5651 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__conb_1_32/HI 7.93e-21
C5652 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -0.00602f
C5653 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# V_LOW 0.0265f
C5654 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# -1.44e-20
C5655 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 4.66e-19
C5656 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.00106f
C5657 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 5.05e-19
C5658 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 0.00122f
C5659 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_12/HI 1.8e-20
C5660 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# -3.57e-19
C5661 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# -3.86e-20
C5662 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0.011f
C5663 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_67/A 0.00479f
C5664 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__conb_1_41/HI 1.58e-19
C5665 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# -3.79e-20
C5666 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# -0.00336f
C5667 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00882f
C5668 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# V_LOW 0.0142f
C5669 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# 0.00216f
C5670 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.24e-21
C5671 sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__conb_1_16/HI 3.35e-19
C5672 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.43e-21
C5673 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_48/Y 1.14e-19
C5674 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# V_LOW 0.0421f
C5675 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 3.65e-19
C5676 sky130_fd_sc_hd__nor2_1_0/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.227f
C5677 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# CLOCK_GEN.SR_Op.Q 4.2e-19
C5678 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 1.13e-19
C5679 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 1.08e-19
C5680 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 0.0072f
C5681 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 0.00589f
C5682 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 3.11e-19
C5683 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 1.93e-19
C5684 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 2.85e-20
C5685 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 2.52e-21
C5686 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 1.53e-21
C5687 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 1.13e-21
C5688 sky130_fd_sc_hd__conb_1_25/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00576f
C5689 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_66/A 0.172f
C5690 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q -2.62e-20
C5691 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__nand2_1_5/Y 0.0107f
C5692 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 1.6e-20
C5693 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_9/A 0.00187f
C5694 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 2.47e-20
C5695 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.76e-19
C5696 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.88e-19
C5697 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0301f
C5698 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_581_47# -7.91e-19
C5699 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# -0.00631f
C5700 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# -0.0109f
C5701 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.63e-20
C5702 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_31/HI -0.0139f
C5703 sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 4.34e-19
C5704 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/Q_N 7.19e-19
C5705 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 5.81e-19
C5706 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 2.72e-20
C5707 FULL_COUNTER.COUNT_SUB_DFF11.Q V_LOW 2.68f
C5708 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# V_LOW 1.22e-20
C5709 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_381_47# -2.53e-20
C5710 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# sky130_fd_sc_hd__conb_1_46/HI -6.57e-19
C5711 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00484f
C5712 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# V_LOW 0.0114f
C5713 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_7/Y 0.023f
C5714 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/Q_N -8.88e-34
C5715 sky130_fd_sc_hd__inv_16_49/A sky130_fd_sc_hd__inv_16_51/Y 0.00539f
C5716 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_66/A 3.68e-20
C5717 sky130_fd_sc_hd__conb_1_5/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 6.53e-21
C5718 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__conb_1_24/HI 4.46e-19
C5719 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__conb_1_28/HI 0.0137f
C5720 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__inv_1_29/Y 0.00148f
C5721 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_381_47# -3.79e-20
C5722 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# -4.66e-20
C5723 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.53e-20
C5724 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_45/Y 4.56e-21
C5725 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 7.23e-19
C5726 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# V_LOW -2.68e-19
C5727 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00235f
C5728 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_35/Y 5.25e-21
C5729 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__inv_1_41/Y 0.0106f
C5730 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_19/HI 0.0446f
C5731 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.61e-19
C5732 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__conb_1_5/HI 0.00344f
C5733 sky130_fd_sc_hd__conb_1_0/LO RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0115f
C5734 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.0036f
C5735 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 9.65e-21
C5736 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.13e-21
C5737 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 5.74e-19
C5738 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 5.82e-20
C5739 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_1_33/Y 0.00113f
C5740 sky130_fd_sc_hd__dfbbn_1_41/Q_N FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.21e-19
C5741 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 7.12e-19
C5742 sky130_fd_sc_hd__conb_1_25/LO FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.43e-20
C5743 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# sky130_fd_sc_hd__inv_1_44/A 6.11e-19
C5744 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0815f
C5745 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# -9.48e-19
C5746 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# sky130_fd_sc_hd__conb_1_32/HI 1.66e-19
C5747 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 0.00539f
C5748 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.0274f
C5749 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# V_LOW -0.00427f
C5750 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 8.84e-20
C5751 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_40/Y 0.0308f
C5752 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 4.17e-20
C5753 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_47/Y 0.00878f
C5754 sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_8/Y 0.00658f
C5755 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# -2.57e-20
C5756 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF14.Q 0.442f
C5757 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_5/A 0.00457f
C5758 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# sky130_fd_sc_hd__conb_1_25/HI 1.25e-21
C5759 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_28/Y 5.94e-20
C5760 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# sky130_fd_sc_hd__inv_1_13/Y 1.19e-20
C5761 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.185f
C5762 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 0.00126f
C5763 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__conb_1_0/HI 0.00244f
C5764 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_1_33/Y 6.73e-20
C5765 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 1.37e-21
C5766 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# V_LOW 6.78e-19
C5767 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__inv_1_10/Y 0.00117f
C5768 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 6.63e-19
C5769 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 1.01e-19
C5770 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.46e-19
C5771 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# V_LOW -1.01e-19
C5772 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__conb_1_21/HI 7.35e-19
C5773 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 1.97e-19
C5774 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_791_47# 5.19e-19
C5775 sky130_fd_sc_hd__inv_16_22/A sky130_fd_sc_hd__inv_16_8/Y 6.16e-19
C5776 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00211f
C5777 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 9.56e-19
C5778 V_SENSE sky130_fd_sc_hd__conb_1_47/HI 7.21e-19
C5779 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0325f
C5780 sky130_fd_sc_hd__conb_1_25/HI FALLING_COUNTER.COUNT_SUB_DFF12.Q 7.24e-19
C5781 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 5.75e-22
C5782 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 4.4e-21
C5783 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__inv_1_64/Y 7.41e-22
C5784 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 9.61e-21
C5785 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.00192f
C5786 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__conb_1_6/HI 0.00139f
C5787 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__inv_16_42/Y 0.0197f
C5788 sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__conb_1_17/HI 0.026f
C5789 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# V_LOW 0.00622f
C5790 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_29/LO 8.81e-20
C5791 V_SENSE sky130_fd_sc_hd__conb_1_44/LO 9.19e-19
C5792 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_49/A 0.0272f
C5793 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# V_LOW 2.26e-20
C5794 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_193_47# 0.318f
C5795 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00112f
C5796 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# 0.0179f
C5797 sky130_fd_sc_hd__nand3_1_1/a_193_47# sky130_fd_sc_hd__nand3_1_1/Y 3.9e-19
C5798 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# sky130_fd_sc_hd__inv_1_69/Y 5.11e-19
C5799 Reset sky130_fd_sc_hd__inv_1_44/A 0.451f
C5800 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_44/A 0.00143f
C5801 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 7.94e-20
C5802 sky130_fd_sc_hd__dfbbn_1_33/Q_N V_LOW -0.00993f
C5803 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_33/HI 0.206f
C5804 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# -1.44e-20
C5805 sky130_fd_sc_hd__inv_1_60/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0582f
C5806 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00173f
C5807 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# V_LOW 4.8e-20
C5808 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_42/Y 5.93e-20
C5809 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 7.91e-20
C5810 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -5.02e-19
C5811 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# -0.00344f
C5812 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# 0.00278f
C5813 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_1_58/Y 0.113f
C5814 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__inv_16_41/Y 1.64e-19
C5815 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__conb_1_28/HI -0.00262f
C5816 RISING_COUNTER.COUNT_SUB_DFF1.Q transmission_gate_9/GN 2.34e-19
C5817 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__inv_1_29/Y 0.0126f
C5818 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_16_4/Y 0.038f
C5819 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__conb_1_45/HI 1.79e-21
C5820 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16_51/A 0.00341f
C5821 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.039f
C5822 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 0.00438f
C5823 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.74e-21
C5824 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__conb_1_32/HI 2.2e-19
C5825 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__conb_1_5/HI -7.5e-19
C5826 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.00732f
C5827 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__conb_1_20/HI 6.53e-20
C5828 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_1_67/A 0.215f
C5829 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_19/HI 2.24e-20
C5830 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 9.71e-19
C5831 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# Reset 0.0196f
C5832 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_8/HI 0.00174f
C5833 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__inv_16_41/Y 3.56e-19
C5834 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__conb_1_23/HI 0.00967f
C5835 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_30/LO 0.0121f
C5836 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 0.0195f
C5837 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# -0.00813f
C5838 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/Q_N -2.17e-19
C5839 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 3.09e-20
C5840 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 0.00202f
C5841 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 1.76e-20
C5842 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nand2_8_8/A 5.58e-20
C5843 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0114f
C5844 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# -5.54e-21
C5845 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 0.00518f
C5846 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0333f
C5847 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 1.43e-19
C5848 sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_15/Y 0.0124f
C5849 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_9/Y 0.0111f
C5850 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_581_47# 4.99e-19
C5851 sky130_fd_sc_hd__conb_1_42/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0222f
C5852 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# sky130_fd_sc_hd__conb_1_0/HI 0.00211f
C5853 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__inv_1_12/Y 0.0308f
C5854 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 6.7e-21
C5855 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__inv_1_31/Y 1.1e-20
C5856 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.29e-20
C5857 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# V_LOW -1.39e-35
C5858 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 1.55e-20
C5859 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00527f
C5860 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 4.83e-20
C5861 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_2_0/A 1.15e-20
C5862 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6e-20
C5863 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI 1.77e-19
C5864 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 9.66e-19
C5865 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 4.2e-20
C5866 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 2.01e-20
C5867 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00415f
C5868 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 7.33e-19
C5869 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00152f
C5870 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_26/HI 0.0732f
C5871 sky130_fd_sc_hd__conb_1_28/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00156f
C5872 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.44e-19
C5873 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__inv_1_10/Y 1.86e-19
C5874 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__conb_1_6/HI 3.65e-19
C5875 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 5.61e-20
C5876 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.81e-20
C5877 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# -3.48e-20
C5878 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_891_329# -2.2e-20
C5879 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_791_47# 9.35e-19
C5880 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/Q_N 3.68e-21
C5881 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 5.84e-19
C5882 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_28/Y 0.0246f
C5883 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__conb_1_14/LO 7.24e-19
C5884 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# 0.00121f
C5885 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_2_0/A 0.0304f
C5886 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__conb_1_7/HI 6.51e-19
C5887 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_1_59/Y 1.2e-19
C5888 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.35e-20
C5889 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_9/LO 7.52e-20
C5890 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# sky130_fd_sc_hd__inv_1_41/Y 5.74e-20
C5891 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_21/Y 0.0618f
C5892 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.49e-21
C5893 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.62e-21
C5894 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# -2.57e-20
C5895 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00401f
C5896 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__inv_1_29/Y 0.0204f
C5897 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_56/Y 0.075f
C5898 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.15e-19
C5899 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# 0.00115f
C5900 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__conb_1_2/HI 1.36e-19
C5901 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__conb_1_5/HI -2.17e-19
C5902 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1_45/HI 3.45e-21
C5903 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# V_LOW -0.106f
C5904 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_4/Y 0.00223f
C5905 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# 5.6e-19
C5906 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 2.97e-19
C5907 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__inv_1_45/Y 5.94e-19
C5908 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 7.36e-21
C5909 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# V_LOW 4.8e-20
C5910 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__conb_1_19/HI 7.2e-21
C5911 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00246f
C5912 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 0.0159f
C5913 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# Reset 0.00145f
C5914 FULL_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.05e-20
C5915 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# CLOCK_GEN.SR_Op.Q 0.00328f
C5916 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# V_LOW 0.00656f
C5917 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__conb_1_23/HI -2.07e-19
C5918 sky130_fd_sc_hd__conb_1_6/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.155f
C5919 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 6e-20
C5920 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__conb_1_30/LO 4.7e-20
C5921 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 9.93e-22
C5922 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__inv_1_1/Y 0.00931f
C5923 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# -0.00107f
C5924 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.18e-19
C5925 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.03f
C5926 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 1.38e-19
C5927 sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_1_67/A 5.07e-19
C5928 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# sky130_fd_sc_hd__inv_1_60/Y 0.00136f
C5929 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# -1.46e-20
C5930 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# -0.00263f
C5931 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF15.Q 9.52e-19
C5932 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.00192f
C5933 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.18e-19
C5934 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# V_LOW 0.0122f
C5935 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__inv_1_14/Y 7.97e-21
C5936 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_1_28/Y 7.35e-20
C5937 sky130_fd_sc_hd__dfbbn_1_25/Q_N V_LOW -2.68e-19
C5938 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.32f
C5939 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.0203f
C5940 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__conb_1_41/HI 0.00105f
C5941 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_40/Y 0.108f
C5942 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# 3.53e-19
C5943 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__conb_1_14/HI 1.76e-21
C5944 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_64/Y 1.42e-19
C5945 Reset sky130_fd_sc_hd__inv_1_64/Y 4.48e-20
C5946 sky130_fd_sc_hd__conb_1_21/LO V_LOW 0.0622f
C5947 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.5e-21
C5948 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__conb_1_4/HI 0.00435f
C5949 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 2.05e-19
C5950 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 5.96e-19
C5951 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__inv_1_38/Y 0.00343f
C5952 sky130_fd_sc_hd__dfbbn_1_26/a_581_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.8e-19
C5953 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.84e-20
C5954 sky130_fd_sc_hd__dfbbn_1_4/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0171f
C5955 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_19/HI 3.08e-19
C5956 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__conb_1_38/HI 0.00432f
C5957 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__conb_1_29/HI 2.87e-19
C5958 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0139f
C5959 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 0.0198f
C5960 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_4/LO 5.36e-20
C5961 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# -5.77e-20
C5962 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# -2.52e-19
C5963 sky130_fd_sc_hd__conb_1_10/LO V_LOW 0.0371f
C5964 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 5.59e-19
C5965 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00109f
C5966 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# -3.46e-20
C5967 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_47/HI 0.011f
C5968 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 3.03e-20
C5969 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 4.68e-21
C5970 sky130_fd_sc_hd__inv_1_34/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00532f
C5971 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_40/Y 0.868f
C5972 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__conb_1_7/HI 8.8e-20
C5973 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 9.49e-20
C5974 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__inv_1_59/Y 2.42e-19
C5975 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_44/A 0.0113f
C5976 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.00458f
C5977 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_891_329# -2.2e-20
C5978 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_19/HI 4.65e-19
C5979 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# -0.00491f
C5980 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_15/HI 1.7e-19
C5981 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# -0.00497f
C5982 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.599f
C5983 sky130_fd_sc_hd__nor2_1_0/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 2.23e-20
C5984 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 6.52e-21
C5985 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__inv_1_55/Y 0.0017f
C5986 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_16_2/Y 3.65e-19
C5987 sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_29/A 4.08e-20
C5988 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_15/HI 0.0842f
C5989 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 1.5e-20
C5990 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_1_43/Y 2.58e-21
C5991 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 1.97e-20
C5992 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 6.26e-20
C5993 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# V_LOW -2.68e-19
C5994 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0016f
C5995 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 5.09e-20
C5996 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 8.79e-22
C5997 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 2.76e-20
C5998 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# V_LOW -0.014f
C5999 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__conb_1_38/HI 0.00551f
C6000 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# -0.00263f
C6001 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1_14/LO 1.07e-19
C6002 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.321f
C6003 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# V_LOW 0.0134f
C6004 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# V_LOW 0.00739f
C6005 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_1_30/Y 6.48e-21
C6006 RISING_COUNTER.COUNT_SUB_DFF2.Q Reset 3.85e-21
C6007 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00544f
C6008 sky130_fd_sc_hd__inv_16_22/A sky130_fd_sc_hd__inv_16_29/A 0.0365f
C6009 sky130_fd_sc_hd__inv_16_15/A sky130_fd_sc_hd__inv_16_28/Y 3.35e-19
C6010 sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF12.Q 3.33e-20
C6011 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/Q_N -4.78e-20
C6012 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# -9.32e-20
C6013 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.111f
C6014 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 3.87e-19
C6015 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# V_LOW -0.32f
C6016 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_37/HI 1.24e-20
C6017 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# V_LOW -9.73e-19
C6018 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# V_LOW 0.00693f
C6019 sky130_fd_sc_hd__dfbbn_1_44/a_557_413# sky130_fd_sc_hd__inv_1_39/Y 8.17e-19
C6020 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0017f
C6021 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_19/HI 0.285f
C6022 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__inv_1_28/Y 1.15e-19
C6023 sky130_fd_sc_hd__conb_1_5/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00111f
C6024 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 1.07e-19
C6025 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 0.00237f
C6026 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_22/A 0.159f
C6027 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 0.0354f
C6028 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__conb_1_41/HI -6.57e-19
C6029 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.3e-19
C6030 sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__inv_16_41/Y 0.428f
C6031 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 0.0278f
C6032 sky130_fd_sc_hd__inv_1_64/A FULL_COUNTER.COUNT_SUB_DFF0.Q 9.59e-20
C6033 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 7.23e-21
C6034 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__inv_1_38/Y 0.00182f
C6035 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00266f
C6036 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_14/Y 0.0021f
C6037 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.66e-20
C6038 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__conb_1_38/HI 0.00138f
C6039 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__conb_1_29/HI 3.29e-20
C6040 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_32/Y 6.8e-19
C6041 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_1_10/Y 6.01e-21
C6042 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__conb_1_26/HI 0.0024f
C6043 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_24/Y 5.9e-19
C6044 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q -3.6e-20
C6045 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# -1.76e-19
C6046 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__conb_1_16/LO 5.58e-20
C6047 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# V_LOW 0.0102f
C6048 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 1.51e-20
C6049 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 0.0113f
C6050 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.13f
C6051 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_25/Y 8.76e-20
C6052 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_29/Y 3.02e-19
C6053 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_47/HI 3.09e-20
C6054 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 6.21e-21
C6055 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 1.07e-19
C6056 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# sky130_fd_sc_hd__conb_1_51/HI 2.11e-19
C6057 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00934f
C6058 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 0.00349f
C6059 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__conb_1_7/HI 7.94e-19
C6060 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 0.206f
C6061 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 8.44e-20
C6062 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# -2.53e-20
C6063 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 0.0107f
C6064 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1_21/Y 0.412f
C6065 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 3.27e-19
C6066 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# sky130_fd_sc_hd__inv_1_44/A 0.00165f
C6067 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__nand2_1_5/Y 0.217f
C6068 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# -1.42e-32
C6069 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# -0.00385f
C6070 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# V_LOW -0.104f
C6071 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0501f
C6072 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__conb_1_6/HI 0.0083f
C6073 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 2.19e-19
C6074 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__conb_1_15/HI 6.53e-19
C6075 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.74e-19
C6076 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.74e-19
C6077 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.99e-20
C6078 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.99e-20
C6079 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.0256f
C6080 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# -1.44e-20
C6081 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.88e-19
C6082 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.57e-19
C6083 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 4.25e-19
C6084 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.156f
C6085 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.76e-21
C6086 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.73e-19
C6087 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__nor2_1_0/Y 0.0296f
C6088 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_891_329# -3.85e-20
C6089 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# -0.00459f
C6090 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 5.96e-21
C6091 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 8.26e-21
C6092 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_27_47# 0.0302f
C6093 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# V_LOW 3.56e-20
C6094 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF17.Q 7.32e-19
C6095 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# V_LOW -0.00585f
C6096 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__inv_1_61/Y 2.78e-20
C6097 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__conb_1_17/HI 1.77e-19
C6098 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# -9.32e-20
C6099 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# V_LOW -0.00389f
C6100 sky130_fd_sc_hd__inv_1_25/Y sky130_fd_sc_hd__inv_16_41/Y 4.66e-19
C6101 sky130_fd_sc_hd__inv_1_38/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00519f
C6102 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__conb_1_29/LO 0.012f
C6103 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00258f
C6104 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# V_LOW 0.00739f
C6105 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0299f
C6106 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 1.03e-19
C6107 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_46/HI 1.88e-19
C6108 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 1.25e-19
C6109 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.38e-19
C6110 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 5.25e-20
C6111 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__conb_1_9/HI 5.87e-20
C6112 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# V_LOW 0.00521f
C6113 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/Q_N -4.33e-20
C6114 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__conb_1_20/HI 0.0632f
C6115 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 5.21e-20
C6116 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 3.01e-21
C6117 sky130_fd_sc_hd__inv_16_8/A V_LOW 0.37f
C6118 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# V_LOW -2.78e-35
C6119 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0325f
C6120 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.0033f
C6121 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.4e-19
C6122 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# 7.63e-19
C6123 sky130_fd_sc_hd__inv_1_23/Y V_LOW 0.159f
C6124 sky130_fd_sc_hd__conb_1_36/HI RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0184f
C6125 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 9.03e-19
C6126 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_16/HI 1.88e-19
C6127 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__inv_1_63/Y 0.00204f
C6128 FALLING_COUNTER.COUNT_SUB_DFF4.Q V_LOW 2.76f
C6129 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 2.51e-19
C6130 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__conb_1_38/HI 1.51e-20
C6131 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 5.96e-19
C6132 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# V_LOW -0.00371f
C6133 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/Q_N 0.00167f
C6134 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_0/Y 0.00123f
C6135 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__conb_1_36/LO 0.00107f
C6136 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_66/A 2.77e-20
C6137 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0397f
C6138 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0262f
C6139 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0122f
C6140 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0244f
C6141 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0357f
C6142 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_48/HI 0.00903f
C6143 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# V_LOW -0.00583f
C6144 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# -1.44e-20
C6145 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 0.00151f
C6146 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 9.67e-20
C6147 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0456f
C6148 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 0.0199f
C6149 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_15/LO 1.13e-21
C6150 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__conb_1_9/HI 0.228f
C6151 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# V_LOW -9.94e-19
C6152 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_647_21# -1.93e-19
C6153 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.00585f
C6154 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# sky130_fd_sc_hd__conb_1_6/HI 5.87e-20
C6155 FALLING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0276f
C6156 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0098f
C6157 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.34e-19
C6158 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_24/LO 1.67e-19
C6159 sky130_fd_sc_hd__inv_16_28/Y sky130_fd_sc_hd__inv_16_8/Y 0.021f
C6160 sky130_fd_sc_hd__inv_16_9/Y sky130_fd_sc_hd__inv_16_8/A 2.72e-19
C6161 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 1.34e-19
C6162 sky130_fd_sc_hd__inv_1_66/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 6.04e-19
C6163 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# V_LOW -0.0165f
C6164 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__inv_1_55/Y 2.81e-19
C6165 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0141f
C6166 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__conb_1_33/HI 1.36e-20
C6167 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 1.11e-20
C6168 sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00105f
C6169 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# sky130_fd_sc_hd__conb_1_8/HI -6.57e-19
C6170 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 1.17e-20
C6171 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 2.18e-19
C6172 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 3.64e-20
C6173 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# -0.00552f
C6174 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# -4.66e-20
C6175 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# -3.79e-20
C6176 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 9.69e-21
C6177 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 2.95e-22
C6178 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 3.84e-21
C6179 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 3.79e-21
C6180 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00168f
C6181 sky130_fd_sc_hd__conb_1_35/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00697f
C6182 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/Q_N -4.24e-20
C6183 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 0.304f
C6184 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0197f
C6185 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_2/Y 0.0035f
C6186 sky130_fd_sc_hd__conb_1_5/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 3.91e-20
C6187 V_SENSE sky130_fd_sc_hd__conb_1_46/LO 9.19e-19
C6188 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# V_LOW 0.0165f
C6189 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 2.82e-19
C6190 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 4.03e-19
C6191 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 0.0116f
C6192 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 0.0116f
C6193 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 0.00278f
C6194 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 0.00114f
C6195 sky130_fd_sc_hd__dfbbn_1_36/Q_N FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0167f
C6196 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_193_47# -0.0152f
C6197 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_557_413# -0.0012f
C6198 sky130_fd_sc_hd__dfbbn_1_2/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.43e-19
C6199 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# -0.0244f
C6200 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 9.45e-20
C6201 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.35e-20
C6202 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# V_LOW -2.78e-35
C6203 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0868f
C6204 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0.0272f
C6205 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0489f
C6206 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__conb_1_37/HI 0.0269f
C6207 sky130_fd_sc_hd__dfbbn_1_29/Q_N V_LOW -0.00509f
C6208 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__conb_1_0/HI 3.6e-19
C6209 FALLING_COUNTER.COUNT_SUB_DFF1.Q Reset 0.358f
C6210 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_29/Y 0.297f
C6211 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0196f
C6212 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 8.86e-19
C6213 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.02e-19
C6214 sky130_fd_sc_hd__nand3_1_1/a_193_47# V_LOW -5.03e-19
C6215 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16_51/Y 2.79e-19
C6216 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_49/A 0.116f
C6217 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 9.76e-19
C6218 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.43e-22
C6219 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0237f
C6220 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_8_0/A 8.68e-20
C6221 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__conb_1_50/HI -0.00294f
C6222 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__conb_1_9/HI 0.0289f
C6223 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# -3.79e-20
C6224 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# -4.66e-20
C6225 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__conb_1_8/HI 4.49e-20
C6226 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 5.59e-20
C6227 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__nand3_1_1/Y 1.51e-19
C6228 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# -7.77e-19
C6229 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# -0.0125f
C6230 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.85e-20
C6231 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 5.88e-19
C6232 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 7.67e-19
C6233 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 0.00863f
C6234 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 1.62e-19
C6235 FULL_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0282f
C6236 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__inv_1_39/Y 6.09e-21
C6237 sky130_fd_sc_hd__conb_1_6/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.447f
C6238 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF18.Q 0.184f
C6239 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_1_22/Y 3.38e-19
C6240 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00477f
C6241 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0183f
C6242 FALLING_COUNTER.COUNT_SUB_DFF2.Q Reset 0.00237f
C6243 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__conb_1_10/HI 1.11e-19
C6244 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_1_5/Y 9.68e-19
C6245 sky130_fd_sc_hd__inv_1_13/Y V_LOW 0.406f
C6246 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__conb_1_48/HI -0.0125f
C6247 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00126f
C6248 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/Q_N 0.0173f
C6249 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 0.00209f
C6250 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 9.12e-21
C6251 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 7.09e-19
C6252 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 2.37e-19
C6253 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.319f
C6254 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 0.00113f
C6255 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__nand3_1_2/Y 2.08e-20
C6256 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__inv_1_59/Y 1.91e-20
C6257 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_31/Y 2.38e-20
C6258 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00136f
C6259 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_1_18/A 5.69e-21
C6260 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 0.0375f
C6261 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 3.75e-20
C6262 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 3.75e-20
C6263 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -0.00864f
C6264 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 0.012f
C6265 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# -6.23e-21
C6266 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -9.88e-20
C6267 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_381_47# -4.37e-20
C6268 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# 5.1e-19
C6269 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_16_2/Y 0.00357f
C6270 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.89e-19
C6271 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# sky130_fd_sc_hd__inv_1_0/Y 5.03e-19
C6272 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# V_LOW -6.55e-19
C6273 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_891_329# -2.2e-20
C6274 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# -0.00198f
C6275 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00985f
C6276 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0313f
C6277 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__inv_1_41/Y 3.44e-19
C6278 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__inv_1_38/Y 0.0277f
C6279 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00142f
C6280 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 3.79e-21
C6281 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 9.79e-21
C6282 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 1.12e-20
C6283 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/Q_N -4.97e-19
C6284 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 3.54e-21
C6285 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 5.18e-21
C6286 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 4.13e-21
C6287 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.42e-19
C6288 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 3.53e-21
C6289 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 1.03e-19
C6290 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 2.75e-20
C6291 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__conb_1_46/HI 2.83e-20
C6292 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.0141f
C6293 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.81e-19
C6294 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# V_LOW 0.0124f
C6295 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00314f
C6296 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_1_46/A 0.0591f
C6297 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0.00122f
C6298 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 5.05e-19
C6299 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.00106f
C6300 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 4.66e-19
C6301 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__conb_1_20/HI 1.67e-19
C6302 sky130_fd_sc_hd__dfbbn_1_46/Q_N V_LOW -0.00152f
C6303 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_16_4/Y 2.41e-19
C6304 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_891_329# 2.21e-20
C6305 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.036f
C6306 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00499f
C6307 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0033f
C6308 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__conb_1_0/HI 1.16e-19
C6309 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__inv_1_47/A 2.83e-20
C6310 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 6.31e-19
C6311 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF9.Q 2.33e-20
C6312 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# 7.02e-20
C6313 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 1.19e-19
C6314 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 6.12e-19
C6315 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 0.00954f
C6316 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__inv_1_26/Y 3.76e-21
C6317 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q -5.45e-20
C6318 sky130_fd_sc_hd__conb_1_41/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.56e-20
C6319 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 4.55e-19
C6320 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 2.99e-21
C6321 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__inv_1_2/Y 0.00163f
C6322 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# V_LOW 0.0143f
C6323 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__inv_1_30/Y 7.86e-20
C6324 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_59/Y 0.00151f
C6325 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_56/A 0.00156f
C6326 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 2.52e-20
C6327 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_891_329# 7.97e-21
C6328 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# -0.00834f
C6329 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -1.61e-19
C6330 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0358f
C6331 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# V_LOW 4.8e-20
C6332 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__conb_1_50/HI -2.07e-19
C6333 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 4.74e-21
C6334 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_2_0/A 3.46e-19
C6335 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__conb_1_3/HI 0.01f
C6336 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# -1.66e-19
C6337 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 3.1e-19
C6338 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 0.00243f
C6339 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_1_9/Y 0.0032f
C6340 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.93e-19
C6341 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__conb_1_30/HI 6.8e-19
C6342 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.05e-20
C6343 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF6.Q 4.07e-20
C6344 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__inv_1_33/Y 9.13e-19
C6345 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0206f
C6346 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__inv_1_40/Y 0.00266f
C6347 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_1_34/Y -2.87e-20
C6348 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00134f
C6349 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 0.014f
C6350 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__conb_1_14/HI 5.21e-19
C6351 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__conb_1_10/HI 2.95e-19
C6352 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__conb_1_27/HI 0.00357f
C6353 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 2.5e-19
C6354 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_9/HI 9.96e-21
C6355 sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0513f
C6356 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_66/A 0.165f
C6357 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__inv_1_63/Y 0.00308f
C6358 sky130_fd_sc_hd__dfbbn_1_42/Q_N FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.031f
C6359 FULL_COUNTER.COUNT_SUB_DFF10.Q V_LOW 1.48f
C6360 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 6.09e-21
C6361 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 6.75e-21
C6362 sky130_fd_sc_hd__inv_1_21/Y V_LOW 0.0778f
C6363 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_27_47# 0.00507f
C6364 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# sky130_fd_sc_hd__inv_1_50/Y 4.09e-19
C6365 sky130_fd_sc_hd__conb_1_5/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 6.2e-20
C6366 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__conb_1_33/HI 6.23e-19
C6367 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 2.48e-20
C6368 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 5.34e-19
C6369 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 5.34e-19
C6370 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# Reset 0.0156f
C6371 sky130_fd_sc_hd__conb_1_7/LO V_LOW 0.0541f
C6372 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# -0.00105f
C6373 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 0.00908f
C6374 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__inv_16_42/Y 0.449f
C6375 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_1_33/Y 1.02e-21
C6376 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.94e-20
C6377 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.61e-19
C6378 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_44/A 0.00207f
C6379 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 5.78e-21
C6380 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__conb_1_7/HI 0.348f
C6381 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1_49/LO 9.25e-19
C6382 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.147f
C6383 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# -0.00385f
C6384 sky130_fd_sc_hd__dfbbn_1_22/Q_N FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0018f
C6385 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__conb_1_2/HI 0.00375f
C6386 sky130_fd_sc_hd__inv_16_40/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0565f
C6387 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_18/LO 0.0541f
C6388 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__inv_1_59/Y 9.37e-19
C6389 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__conb_1_29/HI 7.39e-19
C6390 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.55e-19
C6391 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 1.27e-20
C6392 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 6.86e-21
C6393 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00304f
C6394 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 0.00185f
C6395 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.00411f
C6396 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.58e-20
C6397 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# V_LOW 1.79e-20
C6398 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_1/Y 0.00157f
C6399 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# -0.00117f
C6400 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# -0.00512f
C6401 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_557_413# -0.0012f
C6402 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# -0.00335f
C6403 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# sky130_fd_sc_hd__inv_1_49/Y 1.1e-20
C6404 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00402f
C6405 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# 0.00492f
C6406 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__conb_1_10/HI 1.94e-20
C6407 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0238f
C6408 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00138f
C6409 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_2_0/A 1.09e-20
C6410 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 4.17e-20
C6411 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_3/A 0.181f
C6412 sky130_fd_sc_hd__conb_1_43/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0484f
C6413 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00168f
C6414 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -0.00472f
C6415 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# -2.25e-19
C6416 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_2_0/A 1.28e-19
C6417 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__inv_1_3/Y 0.00318f
C6418 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.21e-19
C6419 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__conb_1_8/LO 8.32e-20
C6420 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.43e-20
C6421 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__inv_1_25/Y 1.04e-19
C6422 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__conb_1_12/HI 5.54e-20
C6423 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00416f
C6424 sky130_fd_sc_hd__inv_1_53/A CLOCK_GEN.SR_Op.Q 5.17e-19
C6425 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# V_LOW 0.0125f
C6426 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# -2.57e-20
C6427 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# -0.00122f
C6428 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# -0.0129f
C6429 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00943f
C6430 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__inv_1_58/Y 0.0977f
C6431 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_1_60/Y 0.0153f
C6432 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 4.16e-19
C6433 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# -3.86e-20
C6434 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_941_21# -5.58e-20
C6435 sky130_fd_sc_hd__inv_1_0/Y Reset 4.89e-20
C6436 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__conb_1_27/HI 0.0247f
C6437 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 3.53e-19
C6438 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_48/Y 1.31e-19
C6439 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.09e-19
C6440 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# V_LOW 1.38e-19
C6441 sky130_fd_sc_hd__inv_1_22/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0927f
C6442 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.039f
C6443 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.208f
C6444 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 8.7e-21
C6445 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 0.0018f
C6446 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.133f
C6447 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_32/LO 5.04e-21
C6448 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 0.00718f
C6449 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__conb_1_9/HI 3.04e-20
C6450 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 8.84e-20
C6451 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00466f
C6452 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.012f
C6453 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 0.375f
C6454 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_1_63/Y 1.43e-19
C6455 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 3.35e-21
C6456 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# 5.75e-19
C6457 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 4.81e-20
C6458 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 9.34e-20
C6459 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 2.04e-19
C6460 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_1_67/A 5.84e-20
C6461 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.44e-20
C6462 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 2.34e-20
C6463 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 6.18e-20
C6464 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_9/Y 0.127f
C6465 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 0.0123f
C6466 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__inv_1_27/Y 1.72e-20
C6467 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# Reset 4.39e-19
C6468 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# sky130_fd_sc_hd__conb_1_23/HI 0.00119f
C6469 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/Q_N -2.17e-19
C6470 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_27/Y 0.0232f
C6471 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# CLOCK_GEN.SR_Op.Q 9.56e-20
C6472 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 3.21e-20
C6473 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 4.41e-21
C6474 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 4.36e-19
C6475 sky130_fd_sc_hd__inv_1_47/A CLOCK_GEN.SR_Op.Q 0.131f
C6476 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/Q_N -6.48e-19
C6477 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_54/Y 0.00171f
C6478 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_66/A 1.98e-21
C6479 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 1.17e-20
C6480 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00275f
C6481 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__conb_1_26/HI 1.97e-19
C6482 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -0.00447f
C6483 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# -2.27e-19
C6484 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_1_26/Y 1.44e-20
C6485 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# -0.00263f
C6486 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -2.18e-19
C6487 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 2.77e-19
C6488 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# -5.54e-21
C6489 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_58/Y 0.321f
C6490 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_25/HI 2.17e-19
C6491 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 0.262f
C6492 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.38e-20
C6493 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# 5.41e-21
C6494 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# 8.79e-22
C6495 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 9.53e-19
C6496 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__inv_1_40/Y 3.02e-21
C6497 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__inv_1_69/Y 1.57e-20
C6498 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.22e-19
C6499 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__nand3_1_2/Y 0.0036f
C6500 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00123f
C6501 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_27/Y 0.0562f
C6502 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 0.00132f
C6503 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0.00113f
C6504 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# -1.64e-19
C6505 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# -7.17e-20
C6506 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# sky130_fd_sc_hd__inv_1_3/Y 1.07e-21
C6507 sky130_fd_sc_hd__conb_1_31/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0183f
C6508 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 0.0125f
C6509 sky130_fd_sc_hd__conb_1_37/HI V_LOW 0.134f
C6510 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 1.86e-20
C6511 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0014f
C6512 sky130_fd_sc_hd__conb_1_46/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00252f
C6513 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.25e-19
C6514 FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.225f
C6515 sky130_fd_sc_hd__inv_1_66/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 6.88e-20
C6516 sky130_fd_sc_hd__conb_1_25/LO FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00468f
C6517 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_66/A 0.104f
C6518 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.00595f
C6519 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 3.12e-19
C6520 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# -0.00472f
C6521 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# -8.23e-19
C6522 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_1_32/Y 4.81e-21
C6523 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# V_LOW -0.00341f
C6524 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# V_LOW 0.00756f
C6525 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.00261f
C6526 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_59/Y 0.0304f
C6527 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# V_LOW -0.0685f
C6528 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_1/a_647_21# 0.0125f
C6529 V_SENSE sky130_fd_sc_hd__inv_16_40/Y 9.28e-21
C6530 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# Reset 0.053f
C6531 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_1_44/A 0.00556f
C6532 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 4.16e-19
C6533 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0.0343f
C6534 sky130_fd_sc_hd__conb_1_35/HI FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0187f
C6535 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# -2.57e-20
C6536 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# V_LOW 0.00606f
C6537 sky130_fd_sc_hd__dfbbn_1_3/Q_N FULL_COUNTER.COUNT_SUB_DFF6.Q 1.07e-19
C6538 FALLING_COUNTER.COUNT_SUB_DFF4.Q V_HIGH 0.297f
C6539 sky130_fd_sc_hd__conb_1_11/HI FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0756f
C6540 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.101f
C6541 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.00684f
C6542 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 0.00269f
C6543 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_38/Y 4.56e-21
C6544 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF19.Q 0.00426f
C6545 sky130_fd_sc_hd__nand2_1_5/Y V_LOW 0.368f
C6546 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# 5.49e-19
C6547 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 7.65e-20
C6548 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 7.65e-20
C6549 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00341f
C6550 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# 0.00152f
C6551 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 3.58e-19
C6552 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00996f
C6553 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__inv_1_29/Y 0.00247f
C6554 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# sky130_fd_sc_hd__inv_1_63/Y 4.08e-19
C6555 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00105f
C6556 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0476f
C6557 sky130_fd_sc_hd__inv_1_46/A FULL_COUNTER.COUNT_SUB_DFF2.Q 1.58e-19
C6558 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 0.292f
C6559 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0381f
C6560 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 3.87e-21
C6561 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.03f
C6562 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 5.37e-20
C6563 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1_32/HI 0.0723f
C6564 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_16_41/Y 2.04e-19
C6565 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# V_LOW 0.0158f
C6566 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 2.29e-20
C6567 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00391f
C6568 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_30/Y 2.48e-19
C6569 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# 0.00206f
C6570 sky130_fd_sc_hd__nand2_8_7/a_27_47# V_LOW -0.0117f
C6571 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_47/A 1.93e-19
C6572 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_67/A 0.0259f
C6573 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 8.6e-19
C6574 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0.0032f
C6575 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.00109f
C6576 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 0.00499f
C6577 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.86e-21
C6578 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0281f
C6579 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# -9.32e-20
C6580 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_13/LO 5.36e-19
C6581 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# -1.66e-19
C6582 sky130_fd_sc_hd__conb_1_6/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00604f
C6583 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__nand2_1_2/A 0.01f
C6584 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__inv_1_32/Y 3.72e-19
C6585 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# V_LOW 2.26e-20
C6586 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__inv_1_28/Y 0.00222f
C6587 sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF14.Q 4.59e-19
C6588 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/Q_N -9.56e-20
C6589 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 6.6e-19
C6590 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# 2.35e-19
C6591 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# 2.04e-19
C6592 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 1.03e-19
C6593 sky130_fd_sc_hd__inv_16_16/Y sky130_fd_sc_hd__inv_16_33/Y 0.0359f
C6594 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_791_47# 4.36e-19
C6595 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 4.3e-19
C6596 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 3.04e-19
C6597 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# 0.00104f
C6598 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_1_36/Y 0.00233f
C6599 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 0.00778f
C6600 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# -0.00263f
C6601 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# -1.46e-20
C6602 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0185f
C6603 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__conb_1_27/LO 0.0131f
C6604 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.03e-19
C6605 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# V_LOW 4.8e-20
C6606 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 0.0058f
C6607 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 0.0113f
C6608 RISING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0264f
C6609 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 5.2e-22
C6610 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 7.8e-20
C6611 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# V_LOW -1.39e-35
C6612 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# V_LOW 0.0146f
C6613 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.011f
C6614 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 3.74e-19
C6615 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_66/Y 1.48e-20
C6616 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.38e-20
C6617 sky130_fd_sc_hd__conb_1_27/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 7.65e-19
C6618 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# V_LOW -2.68e-19
C6619 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00276f
C6620 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# -4.66e-20
C6621 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# -3.79e-20
C6622 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__conb_1_16/HI -0.00234f
C6623 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -0.00932f
C6624 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# -0.012f
C6625 sky130_fd_sc_hd__inv_16_6/A V_LOW 0.814f
C6626 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__inv_1_44/A 6.38e-20
C6627 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_1_7/Y 1.24e-21
C6628 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.77e-20
C6629 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# V_LOW 1.38e-19
C6630 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# sky130_fd_sc_hd__nor2_1_0/Y 4.65e-20
C6631 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_1_24/Y 5.41e-22
C6632 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1_22/LO 0.00126f
C6633 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# -2.14e-19
C6634 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# -2.74e-21
C6635 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# -7.6e-19
C6636 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 0.0127f
C6637 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 4.58e-19
C6638 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 7.44e-21
C6639 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 2.38e-20
C6640 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00122f
C6641 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 6.1e-21
C6642 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__inv_1_43/Y 0.00534f
C6643 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_26/HI 0.188f
C6644 RISING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF2.Q 1.71f
C6645 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.0417f
C6646 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__conb_1_41/HI 1.68e-19
C6647 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# -0.00144f
C6648 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# V_LOW 1.79e-20
C6649 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_39/Y 0.00383f
C6650 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__conb_1_30/HI 0.00267f
C6651 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 9.29e-21
C6652 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__inv_1_30/Y 0.00114f
C6653 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_2/HI 0.151f
C6654 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# sky130_fd_sc_hd__inv_1_8/Y 4.43e-19
C6655 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_8/HI 0.0243f
C6656 sky130_fd_sc_hd__inv_16_4/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0292f
C6657 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.81e-20
C6658 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.018f
C6659 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 3.27e-20
C6660 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_28/LO 2.61e-19
C6661 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 5.84e-20
C6662 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nor2_1_0/Y 2.11e-19
C6663 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# V_LOW 0.0232f
C6664 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 4.61e-19
C6665 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 6.96e-19
C6666 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 4.1e-19
C6667 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__conb_1_8/HI 0.00229f
C6668 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/Q_N -4.78e-20
C6669 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0231f
C6670 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00102f
C6671 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_9/Y 9.57e-22
C6672 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00219f
C6673 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 6.39e-20
C6674 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00286f
C6675 RISING_COUNTER.COUNT_SUB_DFF6.Q V_LOW 2.28f
C6676 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# 1.98e-20
C6677 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# 2.72e-19
C6678 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# V_LOW 4.8e-20
C6679 sky130_fd_sc_hd__inv_1_67/Y V_LOW 0.0728f
C6680 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# -0.0103f
C6681 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# -0.00258f
C6682 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# V_LOW -0.00987f
C6683 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0975f
C6684 sky130_fd_sc_hd__conb_1_5/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 2.07e-20
C6685 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0358f
C6686 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 4.01e-19
C6687 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__inv_1_36/Y 5.96e-19
C6688 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__inv_1_27/Y 2.72e-20
C6689 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 2.2e-19
C6690 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# 2.98e-19
C6691 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0361f
C6692 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# -9.32e-20
C6693 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# -6.23e-21
C6694 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_381_47# -3.04e-19
C6695 sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__inv_1_66/A 7.91e-19
C6696 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__inv_16_41/Y 0.0216f
C6697 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/Q_N -9.56e-20
C6698 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.39e-20
C6699 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.37e-19
C6700 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__inv_1_35/Y 6.13e-21
C6701 sky130_fd_sc_hd__dfbbn_1_5/Q_N V_LOW -0.0104f
C6702 FALLING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 3.48f
C6703 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_51/A 0.00351f
C6704 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_12/HI 6.83e-19
C6705 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.03e-19
C6706 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_6/LO 0.0157f
C6707 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF12.Q 0.213f
C6708 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# V_LOW -0.00121f
C6709 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.47e-20
C6710 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# sky130_fd_sc_hd__conb_1_16/HI -0.00264f
C6711 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# -2.57e-20
C6712 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__inv_16_41/Y 2.66e-19
C6713 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__inv_1_41/Y 0.00178f
C6714 sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 7.22e-20
C6715 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__inv_16_40/Y 1.03e-20
C6716 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__conb_1_5/HI 4.56e-21
C6717 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/Q_N 0.0215f
C6718 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_48/Y 0.00182f
C6719 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__conb_1_8/HI 5.74e-19
C6720 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_24/HI 0.00283f
C6721 sky130_fd_sc_hd__inv_1_62/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00458f
C6722 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 1.25e-20
C6723 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF17.Q 1.15e-20
C6724 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_23/HI 0.0217f
C6725 sky130_fd_sc_hd__nand2_8_3/a_27_47# CLOCK_GEN.SR_Op.Q 3.76e-19
C6726 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 1.21e-19
C6727 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0311f
C6728 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# 1.21e-19
C6729 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__conb_1_40/HI 6.9e-19
C6730 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# -9.32e-20
C6731 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_17/HI -0.00105f
C6732 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 4.02e-20
C6733 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0307f
C6734 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 8e-21
C6735 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_20/Y 0.0355f
C6736 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_53/Y 6.79e-20
C6737 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 0.0109f
C6738 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0308f
C6739 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_193_47# -0.0595f
C6740 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__conb_1_28/HI 3.94e-20
C6741 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# -0.00141f
C6742 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_2_0/A 4.15e-20
C6743 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__conb_1_19/HI 0.00248f
C6744 sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__inv_1_64/Y 2.76e-19
C6745 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00183f
C6746 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 0.00189f
C6747 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00189f
C6748 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00596f
C6749 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 1.75e-19
C6750 sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_47/Y 0.187f
C6751 sky130_fd_sc_hd__conb_1_33/LO FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.34e-20
C6752 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 0.00441f
C6753 sky130_fd_sc_hd__conb_1_22/HI RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0545f
C6754 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16_49/Y 0.393f
C6755 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.125f
C6756 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI -4.47e-19
C6757 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# V_LOW 0.0122f
C6758 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.49e-19
C6759 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__conb_1_15/HI 0.00359f
C6760 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_1_31/Y 0.00279f
C6761 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_16_8/Y 0.025f
C6762 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_24/HI 0.0277f
C6763 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__conb_1_28/HI 0.00102f
C6764 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0115f
C6765 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 9.98e-20
C6766 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 3.4e-20
C6767 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# -9.41e-19
C6768 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0.00132f
C6769 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00113f
C6770 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 7.04e-19
C6771 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0103f
C6772 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.13e-20
C6773 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# sky130_fd_sc_hd__conb_1_47/HI 2.48e-19
C6774 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 4.07e-20
C6775 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 7e-19
C6776 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__conb_1_25/HI 0.0632f
C6777 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/Q_N -4.33e-20
C6778 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__inv_1_62/Y 2.3e-19
C6779 sky130_fd_sc_hd__inv_16_49/A sky130_fd_sc_hd__inv_16_55/Y 0.00365f
C6780 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.01f
C6781 sky130_fd_sc_hd__fill_8_852/VPB V_LOW 0.797f
C6782 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0363f
C6783 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 2.03e-20
C6784 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# V_LOW 0.0021f
C6785 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__conb_1_29/HI 1.88e-19
C6786 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_381_47# -0.00516f
C6787 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__conb_1_4/HI 0.0129f
C6788 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.32e-19
C6789 V_SENSE Reset 24.8f
C6790 sky130_fd_sc_hd__dfbbn_1_6/Q_N V_LOW -0.0104f
C6791 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.0245f
C6792 FALLING_COUNTER.COUNT_SUB_DFF7.Q V_LOW 0.86f
C6793 sky130_fd_sc_hd__inv_16_26/Y V_LOW 0.256f
C6794 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__conb_1_5/HI 5.88e-20
C6795 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__inv_1_58/Y -5.28e-20
C6796 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__inv_1_14/Y 0.00525f
C6797 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_647_21# -0.00115f
C6798 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# -0.00375f
C6799 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.81e-21
C6800 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__inv_1_66/A 9.78e-19
C6801 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_18/HI 0.122f
C6802 sky130_fd_sc_hd__conb_1_2/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 0.122f
C6803 sky130_fd_sc_hd__conb_1_39/LO V_LOW 0.0684f
C6804 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/Q_N -4.24e-20
C6805 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# V_LOW 0.00245f
C6806 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.21e-19
C6807 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0.00987f
C6808 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0.0101f
C6809 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_1_25/Y 9.74e-20
C6810 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# sky130_fd_sc_hd__conb_1_20/HI 1.25e-21
C6811 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 2.5e-20
C6812 sky130_fd_sc_hd__conb_1_31/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00666f
C6813 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_46/A 2.24e-19
C6814 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 2.07e-20
C6815 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# 1.6e-20
C6816 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# V_LOW 0.0152f
C6817 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# 9.54e-19
C6818 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF13.Q 6.71e-21
C6819 FALLING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 1.24e-20
C6820 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_1_33/Y 2.99e-22
C6821 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 4.09e-19
C6822 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# -0.00279f
C6823 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_891_329# -0.00159f
C6824 Reset sky130_fd_sc_hd__inv_16_41/Y 0.338f
C6825 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.158f
C6826 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_16_41/Y 0.0104f
C6827 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 8.81e-20
C6828 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__conb_1_19/HI -2.07e-19
C6829 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__inv_1_34/Y 1.41e-19
C6830 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.051f
C6831 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_43/Y 2.07e-20
C6832 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.00106f
C6833 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 7.96e-20
C6834 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# 2.71e-19
C6835 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 7.08e-19
C6836 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# sky130_fd_sc_hd__inv_1_29/Y 8.82e-20
C6837 FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.103f
C6838 sky130_fd_sc_hd__conb_1_39/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.211f
C6839 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 0.00101f
C6840 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 0.00483f
C6841 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# V_LOW 0.0116f
C6842 sky130_fd_sc_hd__inv_16_5/A V_LOW 0.312f
C6843 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.045f
C6844 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__conb_1_21/HI -2.07e-19
C6845 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# sky130_fd_sc_hd__inv_1_31/Y 1.38e-20
C6846 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00373f
C6847 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_10/Y 1.5e-19
C6848 sky130_fd_sc_hd__conb_1_5/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.296f
C6849 sky130_fd_sc_hd__inv_16_40/Y CLOCK_GEN.SR_Op.Q 0.0327f
C6850 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__conb_1_30/LO 5.04e-21
C6851 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__conb_1_24/HI -0.0119f
C6852 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_51/Y 1.15e-19
C6853 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# sky130_fd_sc_hd__inv_1_38/Y 6.65e-20
C6854 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__inv_1_37/Y 4.43e-21
C6855 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.021f
C6856 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# Reset 0.00533f
C6857 sky130_fd_sc_hd__conb_1_33/HI RISING_COUNTER.COUNT_SUB_DFF1.Q 6.54e-21
C6858 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_10/HI 0.355f
C6859 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 0.0186f
C6860 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# V_LOW 0.00574f
C6861 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 3.04e-19
C6862 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 4.3e-19
C6863 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_791_47# 4.36e-19
C6864 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 2.52e-19
C6865 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 9.75e-19
C6866 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 1.68e-19
C6867 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00128f
C6868 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_9/LO 9.06e-21
C6869 sky130_fd_sc_hd__conb_1_48/LO FALLING_COUNTER.COUNT_SUB_DFF7.Q 9.36e-21
C6870 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 4.87e-19
C6871 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__inv_1_62/Y 1.54e-20
C6872 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.04e-19
C6873 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_39/Y 3.2e-19
C6874 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0161f
C6875 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__inv_1_47/Y 6.13e-21
C6876 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_25/LO 2.01e-19
C6877 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# -0.0109f
C6878 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_647_21# -6.43e-20
C6879 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0342f
C6880 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.18e-19
C6881 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# Reset 0.0348f
C6882 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__nand2_8_4/Y 5.93e-20
C6883 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# -9.52e-20
C6884 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0366f
C6885 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.94e-20
C6886 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# -0.00107f
C6887 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_40/Y 9.87e-21
C6888 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__conb_1_4/HI 2.25e-19
C6889 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__conb_1_37/HI -0.00182f
C6890 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00321f
C6891 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 6.53e-20
C6892 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 6.03e-20
C6893 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# 5.29e-19
C6894 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_49/A 0.0153f
C6895 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# -0.065f
C6896 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__conb_1_16/HI 0.0132f
C6897 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_581_47# -7.91e-19
C6898 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_1_18/A 0.0121f
C6899 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# -0.00141f
C6900 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 8.39e-20
C6901 sky130_fd_sc_hd__inv_1_19/Y sky130_fd_sc_hd__inv_16_2/Y 4.29e-20
C6902 sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0403f
C6903 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 1.61e-19
C6904 sky130_fd_sc_hd__dfbbn_1_49/Q_N RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00969f
C6905 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 3.44e-20
C6906 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0836f
C6907 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 2.65e-20
C6908 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 3e-19
C6909 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# V_LOW 0.013f
C6910 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_18/HI 0.00128f
C6911 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# -3.79e-20
C6912 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# -0.00336f
C6913 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_647_21# 0.00382f
C6914 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__conb_1_14/HI 5.76e-21
C6915 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# -0.00385f
C6916 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 8.74e-20
C6917 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__conb_1_11/HI -1.96e-19
C6918 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.0398f
C6919 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.218f
C6920 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__inv_1_26/Y 2.04e-19
C6921 sky130_fd_sc_hd__nand2_8_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.63e-19
C6922 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# V_LOW -0.0136f
C6923 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# V_LOW 1.79e-20
C6924 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00868f
C6925 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__conb_1_23/HI 0.145f
C6926 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__conb_1_14/LO 1.63e-21
C6927 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 0.00471f
C6928 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.00921f
C6929 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__conb_1_12/HI 0.00306f
C6930 sky130_fd_sc_hd__inv_16_23/A V_LOW 0.0576f
C6931 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0411f
C6932 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_37/Y 8.85e-19
C6933 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_891_329# 1.93e-20
C6934 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00705f
C6935 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__conb_1_11/HI 0.275f
C6936 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_51/Y 2.83e-21
C6937 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.66e-19
C6938 FALLING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 4.49e-21
C6939 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0548f
C6940 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_557_413# -3.67e-20
C6941 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_891_329# -1.42e-19
C6942 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# -5.33e-20
C6943 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# V_LOW -1.39e-35
C6944 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.8e-19
C6945 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0069f
C6946 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.56e-20
C6947 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 4.71e-20
C6948 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 2.01e-20
C6949 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.52e-19
C6950 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00326f
C6951 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00321f
C6952 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_50/HI 0.056f
C6953 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__inv_1_50/Y 0.0709f
C6954 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 2.04e-21
C6955 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 8.65e-19
C6956 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.26f
C6957 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# -0.0637f
C6958 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__inv_1_33/Y 0.0159f
C6959 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# sky130_fd_sc_hd__conb_1_44/HI 0.00119f
C6960 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 8.35e-19
C6961 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0.0336f
C6962 sky130_fd_sc_hd__conb_1_17/LO V_LOW 0.154f
C6963 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__conb_1_16/HI 2.59e-22
C6964 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# sky130_fd_sc_hd__conb_1_43/HI 0.00111f
C6965 sky130_fd_sc_hd__inv_16_4/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0705f
C6966 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_2/Y 1.39e-20
C6967 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# Reset 0.00507f
C6968 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_581_47# -2.6e-20
C6969 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.022f
C6970 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 6.24e-21
C6971 sky130_fd_sc_hd__dfbbn_1_41/Q_N V_LOW 1.99e-19
C6972 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# CLOCK_GEN.SR_Op.Q 2.33e-19
C6973 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__inv_1_28/Y 9.56e-21
C6974 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.251f
C6975 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.1e-21
C6976 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# 2.4e-21
C6977 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 2.6e-19
C6978 sky130_fd_sc_hd__conb_1_28/LO V_LOW 0.141f
C6979 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0395f
C6980 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_193_47# -3.17e-19
C6981 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 2.63e-19
C6982 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_29/LO 5.37e-20
C6983 sky130_fd_sc_hd__inv_16_6/A V_HIGH 0.796f
C6984 sky130_fd_sc_hd__conb_1_39/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 0.173f
C6985 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 5.25e-21
C6986 sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 0.335f
C6987 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.438f
C6988 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__inv_1_36/Y 1.64e-19
C6989 FALLING_COUNTER.COUNT_SUB_DFF5.Q V_LOW 2.58f
C6990 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# -0.0129f
C6991 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# -0.00122f
C6992 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0338f
C6993 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00385f
C6994 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 2.2e-19
C6995 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# 4.17e-19
C6996 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_16/HI 5.64e-19
C6997 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0426f
C6998 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_1_49/Y 3.89e-20
C6999 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 6.42e-21
C7000 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# V_LOW 1.38e-19
C7001 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# -4.1e-19
C7002 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_891_329# -2.2e-20
C7003 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_891_329# 0.00162f
C7004 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__inv_1_38/Y 8.52e-21
C7005 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# V_LOW 1.79e-20
C7006 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_18/A 7.81e-20
C7007 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__conb_1_18/HI 0.00643f
C7008 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# V_LOW 0.00545f
C7009 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0904f
C7010 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0059f
C7011 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_24/A 0.391f
C7012 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_16_29/A 0.0246f
C7013 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__conb_1_5/HI 0.00123f
C7014 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 1.79e-19
C7015 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 2.1e-19
C7016 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# sky130_fd_sc_hd__inv_1_12/Y 2.58e-21
C7017 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_193_47# -0.11f
C7018 sky130_fd_sc_hd__inv_16_16/Y sky130_fd_sc_hd__inv_16_15/Y 0.00132f
C7019 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.33e-19
C7020 sky130_fd_sc_hd__nand2_1_3/a_113_47# CLOCK_GEN.SR_Op.Q 9.11e-20
C7021 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_24/Y 0.00136f
C7022 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# -3.34e-20
C7023 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0176f
C7024 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 4.01e-20
C7025 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# V_LOW 0.00857f
C7026 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 0.00684f
C7027 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__conb_1_11/HI 8.59e-20
C7028 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0859f
C7029 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00469f
C7030 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 2.73e-20
C7031 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.446f
C7032 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_56/A 0.015f
C7033 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# V_LOW 0.00205f
C7034 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_7/A 3.35e-20
C7035 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI 8.58e-19
C7036 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0386f
C7037 sky130_fd_sc_hd__inv_1_37/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.2e-20
C7038 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00274f
C7039 sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16_48/A 0.00727f
C7040 sky130_fd_sc_hd__conb_1_2/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.338f
C7041 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0852f
C7042 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__inv_1_43/Y 0.00179f
C7043 sky130_fd_sc_hd__inv_16_32/Y V_LOW 0.302f
C7044 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_44/A 0.0276f
C7045 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00146f
C7046 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.3e-19
C7047 sky130_fd_sc_hd__inv_1_60/Y V_LOW 0.188f
C7048 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00558f
C7049 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_381_47# 1.22e-20
C7050 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_1_21/Y 3.08e-21
C7051 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# V_LOW 0.00684f
C7052 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 0.0035f
C7053 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.0029f
C7054 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0.00106f
C7055 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 8.02e-20
C7056 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# -7.77e-19
C7057 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# -2.15e-19
C7058 sky130_fd_sc_hd__dfbbn_1_8/Q_N V_LOW -0.00245f
C7059 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 4.74e-20
C7060 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_25/HI 5.58e-21
C7061 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 0.0026f
C7062 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.87e-21
C7063 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 4.57e-20
C7064 sky130_fd_sc_hd__conb_1_50/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.384f
C7065 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 7.83e-19
C7066 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00618f
C7067 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# V_LOW 0.0127f
C7068 sky130_fd_sc_hd__fill_4_188/VPB V_LOW 0.797f
C7069 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 0.00159f
C7070 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 3.19e-20
C7071 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# V_LOW -0.307f
C7072 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 6.18e-20
C7073 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 5.86e-21
C7074 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_23/Y 0.0153f
C7075 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_16_2/Y 1.95e-19
C7076 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 7.14e-20
C7077 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 4.49e-19
C7078 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 5.31e-19
C7079 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 5.82e-20
C7080 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 1.46e-19
C7081 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0467f
C7082 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 0.0029f
C7083 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.69e-21
C7084 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/Q_N 3.07e-20
C7085 sky130_fd_sc_hd__conb_1_18/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 1.8e-20
C7086 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.18e-21
C7087 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# 3.65e-19
C7088 sky130_fd_sc_hd__conb_1_42/HI FALLING_COUNTER.COUNT_SUB_DFF1.Q 7.01e-20
C7089 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00102f
C7090 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_791_47# -0.00686f
C7091 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 6.84e-21
C7092 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_33/HI -0.00443f
C7093 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 0.00348f
C7094 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.2e-19
C7095 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 5.71e-21
C7096 sky130_fd_sc_hd__dfbbn_1_33/a_581_47# sky130_fd_sc_hd__inv_1_36/Y 2.34e-19
C7097 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_47/Y 2.07e-19
C7098 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0299f
C7099 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -0.00408f
C7100 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# -0.0103f
C7101 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.6e-19
C7102 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__conb_1_31/HI -0.00175f
C7103 sky130_fd_sc_hd__inv_16_32/Y sky130_fd_sc_hd__inv_16_9/Y 0.133f
C7104 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 2.29e-19
C7105 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0209f
C7106 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 1.04e-19
C7107 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# -0.00385f
C7108 sky130_fd_sc_hd__inv_16_32/A V_LOW 0.184f
C7109 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_557_413# -3.67e-20
C7110 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# -0.00182f
C7111 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 4.56e-21
C7112 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.65e-19
C7113 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 8.25e-19
C7114 sky130_fd_sc_hd__conb_1_17/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 1.53e-19
C7115 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# V_LOW 0.062f
C7116 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 4.54e-19
C7117 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# sky130_fd_sc_hd__conb_1_5/HI 3.23e-21
C7118 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__inv_1_40/Y 8.59e-22
C7119 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.0245f
C7120 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__conb_1_24/HI 3.09e-19
C7121 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nand2_8_8/A 4.63e-19
C7122 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_28/HI 0.00422f
C7123 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.67e-21
C7124 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF14.Q 0.022f
C7125 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 5.81e-19
C7126 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# V_LOW -6.26e-19
C7127 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0297f
C7128 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_1_3/Y 6.55e-20
C7129 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__conb_1_32/HI 1.56e-19
C7130 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_47/Y 0.00635f
C7131 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_9/A 0.076f
C7132 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_16_41/Y 0.179f
C7133 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.00445f
C7134 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.0113f
C7135 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.27e-20
C7136 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 8.77e-20
C7137 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.00174f
C7138 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_33/Y 0.00407f
C7139 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 8.37e-20
C7140 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_20/HI 0.0146f
C7141 sky130_fd_sc_hd__nand2_8_4/Y CLOCK_GEN.SR_Op.Q 0.0929f
C7142 Reset CLOCK_GEN.SR_Op.Q 0.919f
C7143 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__inv_1_44/A 0.00688f
C7144 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__conb_1_23/HI 0.004f
C7145 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_65/A 4.41e-20
C7146 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 0.304f
C7147 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 8.34e-20
C7148 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# -5.92e-19
C7149 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 0.0117f
C7150 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# V_LOW -2.78e-35
C7151 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 5.74e-20
C7152 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# -1.66e-19
C7153 sky130_fd_sc_hd__conb_1_31/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00582f
C7154 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# sky130_fd_sc_hd__inv_1_13/Y 4.45e-20
C7155 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 4.02e-19
C7156 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.6e-20
C7157 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 0.23f
C7158 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 0.00716f
C7159 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__conb_1_0/HI 0.0429f
C7160 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_1_33/Y 2.47e-20
C7161 sky130_fd_sc_hd__inv_1_34/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.2f
C7162 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_21/HI 8.44e-22
C7163 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# V_LOW 1.38e-19
C7164 sky130_fd_sc_hd__conb_1_46/LO FALLING_COUNTER.COUNT_SUB_DFF4.Q 3.81e-20
C7165 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.38e-20
C7166 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_23/HI 0.742f
C7167 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__inv_1_10/Y 4.08e-19
C7168 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.12e-19
C7169 sky130_fd_sc_hd__inv_1_56/Y V_LOW 0.217f
C7170 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_1_45/Y 6.67e-22
C7171 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 7.17e-20
C7172 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.65e-19
C7173 V_SENSE RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00615f
C7174 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/Q_N 1.15e-19
C7175 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_791_47# 4.01e-20
C7176 sky130_fd_sc_hd__fill_4_182/VPB V_LOW 0.797f
C7177 sky130_fd_sc_hd__inv_1_57/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.04e-19
C7178 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 5.71e-19
C7179 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0441f
C7180 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 1.51e-21
C7181 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__inv_1_3/Y 5.82e-19
C7182 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 2.07e-20
C7183 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__conb_1_6/HI 0.0037f
C7184 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 4.74e-20
C7185 sky130_fd_sc_hd__conb_1_5/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.18f
C7186 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# V_LOW -0.0426f
C7187 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# V_LOW 4.8e-20
C7188 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_647_21# 0.0383f
C7189 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.3e-19
C7190 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# -9.41e-19
C7191 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 1.56e-19
C7192 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# sky130_fd_sc_hd__conb_1_31/HI -0.0127f
C7193 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# sky130_fd_sc_hd__inv_1_69/Y 7.97e-21
C7194 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_11/LO 0.0141f
C7195 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 5.13e-19
C7196 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_2/HI 0.00998f
C7197 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# -5.42e-19
C7198 sky130_fd_sc_hd__dfbbn_1_21/Q_N V_LOW 1.99e-19
C7199 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.04e-20
C7200 sky130_fd_sc_hd__inv_16_41/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 0.178f
C7201 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# V_LOW 2.94e-20
C7202 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 9.4e-20
C7203 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -1.89e-19
C7204 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# -3.87e-19
C7205 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# 3.78e-19
C7206 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_5/Y 0.0354f
C7207 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 4.56e-21
C7208 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.74e-19
C7209 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__inv_1_25/Y 4.71e-20
C7210 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_557_413# 9.02e-19
C7211 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0334f
C7212 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00357f
C7213 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00702f
C7214 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 3.53e-19
C7215 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_33/LO 0.02f
C7216 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1_19/LO 0.00331f
C7217 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_41/Y 0.432f
C7218 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_16_2/Y 0.0232f
C7219 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# sky130_fd_sc_hd__conb_1_5/HI -6.57e-19
C7220 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 3.45e-20
C7221 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00269f
C7222 sky130_fd_sc_hd__conb_1_6/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0191f
C7223 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__inv_1_33/Y 0.0212f
C7224 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__conb_1_47/LO 8.84e-20
C7225 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.00239f
C7226 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# V_LOW 0.00346f
C7227 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__conb_1_19/HI 2.13e-21
C7228 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# Reset 0.0633f
C7229 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI 0.0014f
C7230 sky130_fd_sc_hd__dfbbn_1_49/Q_N FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0382f
C7231 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 7.72e-20
C7232 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_47/a_381_47# 1.06e-20
C7233 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_557_413# -0.0012f
C7234 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# -0.00938f
C7235 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 0.00692f
C7236 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00846f
C7237 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 7.35e-20
C7238 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 0.00226f
C7239 sky130_fd_sc_hd__dfbbn_1_38/Q_N V_LOW -2.68e-19
C7240 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# -0.00117f
C7241 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# -0.00538f
C7242 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0212f
C7243 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 0.00286f
C7244 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# sky130_fd_sc_hd__conb_1_0/HI 4.8e-19
C7245 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0262f
C7246 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__inv_1_31/Y 0.0133f
C7247 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 4.78e-21
C7248 sky130_fd_sc_hd__conb_1_19/LO RISING_COUNTER.COUNT_SUB_DFF15.Q 2.39e-20
C7249 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.19e-20
C7250 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.9e-19
C7251 V_SENSE sky130_fd_sc_hd__inv_1_62/Y 5.81e-19
C7252 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0103f
C7253 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00321f
C7254 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# sky130_fd_sc_hd__conb_1_11/HI 6.22e-22
C7255 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 9.82e-19
C7256 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 1.71e-19
C7257 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.0015f
C7258 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 1.01e-19
C7259 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0126f
C7260 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__conb_1_14/HI 4.83e-19
C7261 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00152f
C7262 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00102f
C7263 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__inv_1_10/Y 3.86e-19
C7264 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# V_LOW -2.68e-19
C7265 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 7.34e-20
C7266 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0.00131f
C7267 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 6.3e-19
C7268 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# -4.66e-20
C7269 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 3.14e-19
C7270 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__inv_1_28/Y 0.0714f
C7271 sky130_fd_sc_hd__inv_1_4/Y FULL_COUNTER.COUNT_SUB_DFF6.Q 9.04e-20
C7272 FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 5.81f
C7273 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_2_0/A 0.0151f
C7274 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# 4.48e-19
C7275 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0101f
C7276 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 0.121f
C7277 sky130_fd_sc_hd__inv_1_44/A CLOCK_GEN.SR_Op.Q 0.00168f
C7278 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.94e-21
C7279 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__inv_16_40/Y 0.00321f
C7280 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_21/Y 0.00294f
C7281 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# -1.76e-19
C7282 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_2_0/A 1.08e-20
C7283 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 1.55e-20
C7284 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 6.33e-20
C7285 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 3.76e-20
C7286 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00361f
C7287 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.08e-20
C7288 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16_55/Y 0.241f
C7289 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_51/Y 1f
C7290 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 2.51e-20
C7291 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_4_0/A 0.00103f
C7292 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__conb_1_2/HI 4.47e-19
C7293 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# V_LOW 0.00725f
C7294 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__inv_1_1/Y 0.00488f
C7295 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# sky130_fd_sc_hd__inv_16_42/Y 2.39e-20
C7296 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 5.13e-21
C7297 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 9.67e-21
C7298 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 3.51e-20
C7299 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 1.26e-19
C7300 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 0.00124f
C7301 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# V_LOW 2.94e-20
C7302 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 4.68e-21
C7303 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# Reset 6.9e-19
C7304 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.61e-20
C7305 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_46/A 0.0271f
C7306 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# CLOCK_GEN.SR_Op.Q 6.3e-20
C7307 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# V_LOW 0.0112f
C7308 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_21/HI 0.00335f
C7309 sky130_fd_sc_hd__inv_1_10/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0196f
C7310 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__conb_1_23/HI -8.49e-19
C7311 RISING_COUNTER.COUNT_SUB_DFF5.Q V_LOW 1.98f
C7312 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_17/HI 7.44e-22
C7313 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__inv_1_1/Y 5.11e-19
C7314 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_66/A 0.0225f
C7315 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.166f
C7316 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/Q_N 0.00275f
C7317 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 3.68e-19
C7318 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 2.21e-19
C7319 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# sky130_fd_sc_hd__inv_1_60/Y 5.9e-19
C7320 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# -0.00125f
C7321 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# -4.5e-20
C7322 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00196f
C7323 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.335f
C7324 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 7.4e-20
C7325 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# V_LOW 0.00315f
C7326 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_48/Y 2.54e-19
C7327 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__inv_1_14/Y 3.75e-21
C7328 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.0138f
C7329 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.123f
C7330 sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__inv_1_10/Y 2.48e-20
C7331 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_1_19/A 1.62e-19
C7332 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_47/Y 8.12e-19
C7333 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__conb_1_4/HI 0.00255f
C7334 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 2.08e-19
C7335 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_1_38/Y 0.0266f
C7336 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.2e-19
C7337 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__conb_1_14/HI 4.9e-19
C7338 sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 5.59e-20
C7339 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__conb_1_29/HI 0.0132f
C7340 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00435f
C7341 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.627f
C7342 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__conb_1_26/HI 0.00244f
C7343 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# -5.54e-21
C7344 FULL_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0366f
C7345 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_791_47# 4.22e-20
C7346 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__conb_1_47/HI 0.0174f
C7347 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 1.25e-19
C7348 sky130_fd_sc_hd__inv_1_66/A sky130_fd_sc_hd__inv_1_64/A 1.12e-19
C7349 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__inv_2_0/A 0.00199f
C7350 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 1.93e-19
C7351 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_1_46/A 0.445f
C7352 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_44/HI 7.25e-20
C7353 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.26e-20
C7354 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_44/A 0.00157f
C7355 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 3.19e-19
C7356 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# -4.66e-20
C7357 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00894f
C7358 sky130_fd_sc_hd__conb_1_44/LO FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0484f
C7359 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__conb_1_15/HI 5.72e-19
C7360 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_1_21/Y 0.0357f
C7361 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0304f
C7362 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0025f
C7363 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_891_329# -2.46e-19
C7364 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# -0.00717f
C7365 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_557_413# -3.67e-20
C7366 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 3.32e-20
C7367 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 9.26e-21
C7368 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 1.25e-19
C7369 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 7.57e-20
C7370 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__inv_1_55/Y 0.00211f
C7371 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_33/Y 8.06e-21
C7372 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__conb_1_22/LO 8.84e-20
C7373 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_15/HI 0.025f
C7374 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1_14/HI 7.84e-20
C7375 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_1_43/Y 1.14e-21
C7376 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0162f
C7377 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_24/A 7.22e-20
C7378 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# V_LOW -0.00346f
C7379 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.33e-19
C7380 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 6.21e-21
C7381 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_39/Q_N 0.00105f
C7382 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.49e-21
C7383 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# V_LOW -0.00381f
C7384 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_30/Y 0.00118f
C7385 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_52/A 0.243f
C7386 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# CLOCK_GEN.SR_Op.Q 4.98e-19
C7387 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# -0.00125f
C7388 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# -0.00832f
C7389 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# -1.42e-32
C7390 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# V_LOW 1.79e-20
C7391 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__conb_1_23/HI -2.17e-19
C7392 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.13f
C7393 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_41/Y 0.0199f
C7394 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# V_LOW 0.00174f
C7395 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# V_LOW 0.00564f
C7396 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_1_30/Y 2.4e-21
C7397 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00236f
C7398 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.43e-20
C7399 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00235f
C7400 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_67/A 0.295f
C7401 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0468f
C7402 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_37/HI 1.92e-19
C7403 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# V_LOW 0.00852f
C7404 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# V_LOW -0.00387f
C7405 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# sky130_fd_sc_hd__inv_1_39/Y 6.81e-19
C7406 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.85e-19
C7407 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__conb_1_37/HI 2.32e-19
C7408 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_56/A 0.234f
C7409 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__conb_1_39/HI 1.5e-19
C7410 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# sky130_fd_sc_hd__inv_16_40/Y 0.00181f
C7411 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0435f
C7412 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00434f
C7413 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 8.76e-20
C7414 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 0.0171f
C7415 sky130_fd_sc_hd__conb_1_48/HI RISING_COUNTER.COUNT_SUB_DFF10.Q 5.81e-20
C7416 sky130_fd_sc_hd__inv_1_64/Y CLOCK_GEN.SR_Op.Q 0.00142f
C7417 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# sky130_fd_sc_hd__conb_1_4/HI 7.25e-22
C7418 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_31/Y 0.0436f
C7419 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_41/Y 0.0287f
C7420 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_53/A 4.6e-19
C7421 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 2.26e-20
C7422 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 9.59e-20
C7423 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_14/Y 2.9e-19
C7424 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 1.8e-19
C7425 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__conb_1_4/HI 3.21e-21
C7426 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.89e-20
C7427 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# sky130_fd_sc_hd__conb_1_26/HI 0.00215f
C7428 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# -3.34e-20
C7429 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_48/Y 0.0174f
C7430 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# V_LOW 0.00626f
C7431 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_16_41/Y 0.125f
C7432 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_31/Y 7.39e-21
C7433 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_11/LO 0.00601f
C7434 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__inv_1_32/Y 0.00864f
C7435 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.06e-21
C7436 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1_0/Y 0.00267f
C7437 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__conb_1_47/HI 1.73e-19
C7438 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 8.61e-19
C7439 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__conb_1_44/HI 0.00306f
C7440 sky130_fd_sc_hd__inv_16_40/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0289f
C7441 sky130_fd_sc_hd__inv_16_23/Y V_LOW 0.147f
C7442 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# -6.29e-19
C7443 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_557_413# -3.67e-20
C7444 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand2_1_5/Y 0.00557f
C7445 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 5.82e-20
C7446 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_1_59/Y 4.05e-20
C7447 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 9.74e-20
C7448 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.0198f
C7449 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00694f
C7450 RISING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 5.78e-21
C7451 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# V_LOW -0.0144f
C7452 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0411f
C7453 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_16_4/Y 0.0178f
C7454 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 3.06e-19
C7455 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.51e-20
C7456 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 8.15e-20
C7457 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 8.15e-20
C7458 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.51e-20
C7459 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00154f
C7460 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.71e-19
C7461 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 2.6e-19
C7462 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00776f
C7463 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.134f
C7464 sky130_fd_sc_hd__inv_16_3/A V_LOW 0.594f
C7465 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_66/A 0.0888f
C7466 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__conb_1_15/HI 5.26e-20
C7467 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 6.7e-19
C7468 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__conb_1_25/LO 8.81e-20
C7469 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# -0.2f
C7470 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0.0309f
C7471 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# -4.66e-20
C7472 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# -3.79e-20
C7473 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 8.29e-21
C7474 sky130_fd_sc_hd__conb_1_5/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.136f
C7475 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# V_LOW 2.26e-20
C7476 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_193_47# 0.00651f
C7477 RISING_COUNTER.COUNT_SUB_DFF9.Q V_LOW 1.78f
C7478 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q -5.45e-20
C7479 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# V_LOW -1.39e-35
C7480 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 4.92e-21
C7481 sky130_fd_sc_hd__dfbbn_1_43/a_557_413# V_LOW -9.15e-19
C7482 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__conb_1_29/LO 0.00229f
C7483 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0623f
C7484 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__conb_1_16/HI 0.00115f
C7485 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# V_LOW -1.39e-35
C7486 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 7.94e-20
C7487 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 5.92e-19
C7488 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.74e-19
C7489 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.72e-19
C7490 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# V_LOW 1.38e-19
C7491 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__conb_1_20/HI 0.0438f
C7492 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/Q_N -9.56e-20
C7493 RISING_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00309f
C7494 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 0.00228f
C7495 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0512f
C7496 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__conb_1_37/HI 3.29e-20
C7497 sky130_fd_sc_hd__inv_1_12/Y V_LOW 0.0825f
C7498 sky130_fd_sc_hd__dfbbn_1_17/Q_N V_LOW -0.00493f
C7499 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__inv_1_28/Y 1.51e-20
C7500 FALLING_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.08f
C7501 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0299f
C7502 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 1.3e-19
C7503 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__inv_1_1/Y 1.6e-19
C7504 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.21e-19
C7505 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00224f
C7506 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__inv_1_13/Y 0.0014f
C7507 sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF9.Q 2.95e-20
C7508 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# -0.189f
C7509 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_381_47# 0.0211f
C7510 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 4.12e-19
C7511 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# V_LOW -9.15e-19
C7512 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/Q_N -4.78e-20
C7513 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_47/A 7.13e-21
C7514 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__conb_1_36/LO 0.0121f
C7515 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__conb_1_47/HI 6.66e-20
C7516 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00266f
C7517 sky130_fd_sc_hd__inv_1_22/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.278f
C7518 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0823f
C7519 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.6e-19
C7520 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0168f
C7521 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# V_LOW -0.122f
C7522 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__conb_1_48/HI 0.00208f
C7523 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# 3.78e-20
C7524 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0294f
C7525 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.4e-19
C7526 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_53/A 3.79e-19
C7527 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.00335f
C7528 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_15/LO 3.28e-20
C7529 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# V_LOW -0.00333f
C7530 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0416f
C7531 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_473_413# -6.12e-19
C7532 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_48/LO 0.00198f
C7533 sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# sky130_fd_sc_hd__conb_1_6/HI 1.61e-19
C7534 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 9.67e-20
C7535 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.179f
C7536 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0197f
C7537 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 0.0371f
C7538 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 2.56e-19
C7539 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 2.56e-19
C7540 sky130_fd_sc_hd__nand2_1_2/A V_LOW 0.142f
C7541 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_16_40/Y 0.285f
C7542 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_15/LO 0.00154f
C7543 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.0392f
C7544 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# V_LOW -0.327f
C7545 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 3.48e-20
C7546 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_50/LO 1.18e-20
C7547 sky130_fd_sc_hd__conb_1_4/LO V_LOW 0.0454f
C7548 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 0.00153f
C7549 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_19/A 0.172f
C7550 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# 9.52e-19
C7551 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 4.97e-20
C7552 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_791_47# 9.14e-19
C7553 sky130_fd_sc_hd__dfbbn_1_42/Q_N V_LOW -0.0104f
C7554 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/Q_N -9.56e-20
C7555 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00399f
C7556 FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF0.Q 2.74f
C7557 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# V_LOW 0.0113f
C7558 sky130_fd_sc_hd__dfbbn_1_3/Q_N V_LOW -9.29e-19
C7559 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 5.18e-20
C7560 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 1e-19
C7561 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 9.14e-19
C7562 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 7.34e-19
C7563 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_647_21# -0.00149f
C7564 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_21/HI 4.57e-19
C7565 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_891_329# -0.00159f
C7566 sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.97e-19
C7567 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# -0.00882f
C7568 sky130_fd_sc_hd__inv_1_30/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0405f
C7569 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 4.89e-20
C7570 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF17.Q 5.72e-21
C7571 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__conb_1_20/HI 0.0183f
C7572 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 6.17e-20
C7573 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 6.17e-20
C7574 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 1.74e-19
C7575 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.74e-19
C7576 sky130_fd_sc_hd__inv_1_59/Y sky130_fd_sc_hd__inv_1_58/Y 4.59e-20
C7577 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_47/A 0.0161f
C7578 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0354f
C7579 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0205f
C7580 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_64/A 1.19e-20
C7581 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__conb_1_0/HI 1.23e-19
C7582 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_1_47/A 9.36e-21
C7583 sky130_fd_sc_hd__inv_1_60/Y sky130_fd_sc_hd__conb_1_47/HI 5.18e-19
C7584 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_46/LO 6.15e-19
C7585 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__conb_1_14/HI 0.00338f
C7586 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0199f
C7587 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# sky130_fd_sc_hd__conb_1_24/HI 0.00119f
C7588 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 4.97e-20
C7589 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 8.51e-20
C7590 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__conb_1_15/HI 0.00283f
C7591 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0015f
C7592 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0124f
C7593 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# V_LOW 0.058f
C7594 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__conb_1_50/HI -0.00961f
C7595 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0142f
C7596 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_16_4/Y 3.72e-19
C7597 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__conb_1_9/HI 0.0229f
C7598 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_50/Y 0.00281f
C7599 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# -0.00226f
C7600 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# -7.6e-19
C7601 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.01e-19
C7602 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00378f
C7603 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0273f
C7604 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 2.86e-19
C7605 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00174f
C7606 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__inv_1_39/Y 4.43e-21
C7607 sky130_fd_sc_hd__inv_1_10/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0242f
C7608 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# sky130_fd_sc_hd__conb_1_36/LO 4.7e-20
C7609 FULL_COUNTER.COUNT_SUB_DFF9.Q V_LOW 3.35f
C7610 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.38e-19
C7611 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__conb_1_10/HI 2.45e-19
C7612 sky130_fd_sc_hd__dfbbn_1_17/Q_N RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00559f
C7613 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# V_LOW -9.94e-19
C7614 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.166f
C7615 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 7.36e-21
C7616 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.92e-20
C7617 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 4.42e-19
C7618 sky130_fd_sc_hd__inv_1_32/Y FALLING_COUNTER.COUNT_SUB_DFF12.Q 7.09e-19
C7619 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.051f
C7620 V_SENSE sky130_fd_sc_hd__inv_16_48/Y 1.25f
C7621 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 0.403f
C7622 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 5.51e-20
C7623 sky130_fd_sc_hd__inv_1_46/A FULL_COUNTER.COUNT_SUB_DFF1.Q 1.33e-19
C7624 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00954f
C7625 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# -0.00255f
C7626 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__conb_1_43/HI 0.199f
C7627 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_1_31/Y 8.23e-21
C7628 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 3.13e-19
C7629 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_32/Y 4.97e-20
C7630 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 1.05e-19
C7631 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 1.05e-19
C7632 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 5.65e-19
C7633 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_29/Y 0.0202f
C7634 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 2.46e-19
C7635 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_381_47# -2.53e-20
C7636 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 0.277f
C7637 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_67/A 3.54e-19
C7638 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# 7.43e-20
C7639 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# sky130_fd_sc_hd__inv_1_0/Y 0.00162f
C7640 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 9.71e-19
C7641 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_16_40/Y 5.21e-21
C7642 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_1_3/Y 4.55e-20
C7643 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.91e-19
C7644 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# -3.79e-20
C7645 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# -4.66e-20
C7646 RISING_COUNTER.COUNT_SUB_DFF1.Q V_LOW 0.676f
C7647 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/Q_N 8.96e-21
C7648 RISING_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 0.207f
C7649 sky130_fd_sc_hd__conb_1_50/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.2e-19
C7650 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 6.76e-19
C7651 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 8.61e-21
C7652 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 2.1e-21
C7653 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_16/LO 1.7e-20
C7654 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 6.23e-21
C7655 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__inv_16_40/Y 0.041f
C7656 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__inv_16_41/Y 2.84e-20
C7657 RISING_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 9.15e-21
C7658 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.85e-20
C7659 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.0398f
C7660 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_381_47# 1.72e-19
C7661 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00172f
C7662 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# V_LOW 0.0247f
C7663 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_1_49/Y 0.205f
C7664 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0.0298f
C7665 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_581_47# -2.6e-20
C7666 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0272f
C7667 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# -0.00385f
C7668 V_HIGH RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00111f
C7669 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.00106f
C7670 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.0029f
C7671 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0.0035f
C7672 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# 0.00114f
C7673 sky130_fd_sc_hd__inv_1_24/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 7.21e-20
C7674 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.77e-19
C7675 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_16_41/Y 0.594f
C7676 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_64/A 5.61e-21
C7677 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 3.7e-19
C7678 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 0.00315f
C7679 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# 4.44e-19
C7680 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 8.25e-19
C7681 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.48e-22
C7682 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.338f
C7683 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__inv_1_2/Y 0.00466f
C7684 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# V_LOW 0.00904f
C7685 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__inv_1_30/Y 6.22e-19
C7686 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 3.13e-20
C7687 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# sky130_fd_sc_hd__inv_16_41/Y 1.9e-20
C7688 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__conb_1_27/HI 0.00208f
C7689 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# 3.75e-21
C7690 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# -2.35e-19
C7691 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -4.39e-19
C7692 sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# V_LOW 2.94e-20
C7693 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__conb_1_50/HI -0.00166f
C7694 sky130_fd_sc_hd__dfbbn_1_48/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00191f
C7695 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_31/Y 0.021f
C7696 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# sky130_fd_sc_hd__conb_1_9/HI -5.42e-19
C7697 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 7.06e-21
C7698 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.03e-19
C7699 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_1_49/Y 1.94e-22
C7700 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__conb_1_3/HI 0.0188f
C7701 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 0.00196f
C7702 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.44e-19
C7703 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0704f
C7704 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__conb_1_19/HI 0.00119f
C7705 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00511f
C7706 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 8.02e-21
C7707 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00306f
C7708 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_1_34/Y 1.07e-21
C7709 sky130_fd_sc_hd__dfbbn_1_1/Q_N FULL_COUNTER.COUNT_SUB_DFF7.Q 0.018f
C7710 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 0.0398f
C7711 sky130_fd_sc_hd__conb_1_26/LO FALLING_COUNTER.COUNT_SUB_DFF13.Q 3.97e-19
C7712 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# sky130_fd_sc_hd__conb_1_14/HI 9.76e-19
C7713 sky130_fd_sc_hd__conb_1_45/LO sky130_fd_sc_hd__inv_1_61/Y 0.116f
C7714 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 2.04e-19
C7715 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_9/HI 1.17e-21
C7716 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 2.88e-20
C7717 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_1_63/Y 1.13e-19
C7718 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 2.03e-21
C7719 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_193_47# 0.00287f
C7720 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_1_33/Y 0.0272f
C7721 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_791_47# 5.77e-20
C7722 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.392f
C7723 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00856f
C7724 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# sky130_fd_sc_hd__inv_1_50/Y 4.29e-21
C7725 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__conb_1_33/HI 0.00924f
C7726 sky130_fd_sc_hd__inv_16_29/Y sky130_fd_sc_hd__inv_16_22/A 0.13f
C7727 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 3.76e-20
C7728 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# Reset 0.0204f
C7729 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# -6.57e-19
C7730 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 9.13e-21
C7731 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.15f
C7732 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# -1.44e-20
C7733 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__inv_1_33/Y 7.55e-21
C7734 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.3e-19
C7735 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.74e-20
C7736 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00641f
C7737 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__inv_1_3/Y 4.73e-20
C7738 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__conb_1_2/HI 0.00178f
C7739 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__conb_1_33/LO 1.29e-19
C7740 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# sky130_fd_sc_hd__inv_1_59/Y 5.03e-19
C7741 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__conb_1_29/HI 2.06e-20
C7742 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.3e-19
C7743 FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.07e-20
C7744 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.19e-21
C7745 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00169f
C7746 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00487f
C7747 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0.0085f
C7748 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# V_LOW 0.00492f
C7749 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.29e-22
C7750 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# -0.00813f
C7751 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__inv_1_1/Y 0.0046f
C7752 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_891_329# -0.00159f
C7753 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -0.00486f
C7754 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.46e-19
C7755 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 4.68e-21
C7756 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00726f
C7757 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# 5.22e-19
C7758 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__inv_1_40/Y 0.047f
C7759 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_24/HI 0.0369f
C7760 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_5/a_113_47# 2.12e-19
C7761 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 5.74e-20
C7762 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_48/Y 0.0015f
C7763 RISING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF15.Q 2.22f
C7764 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0273f
C7765 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# -0.00138f
C7766 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -7.6e-19
C7767 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_2_0/A 1.94e-20
C7768 sky130_fd_sc_hd__dfbbn_1_34/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0256f
C7769 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__inv_1_3/Y 1.55e-20
C7770 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__conb_1_28/HI 0.0062f
C7771 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__inv_1_2/Y 0.0021f
C7772 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_21/Y 0.00622f
C7773 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__conb_1_51/HI 2.13e-19
C7774 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_5/LO 9.89e-21
C7775 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_51/Y 0.0023f
C7776 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 8.41e-22
C7777 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 9.89e-21
C7778 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/Q_N 2.8e-20
C7779 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_1_25/Y 7.08e-19
C7780 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.00109f
C7781 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# V_LOW 0.00683f
C7782 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# -0.00834f
C7783 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -1.61e-19
C7784 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# -1.66e-19
C7785 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# -7.17e-20
C7786 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00468f
C7787 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_37/HI 0.495f
C7788 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__conb_1_50/HI -2.17e-19
C7789 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.28e-19
C7790 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.09e-19
C7791 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00238f
C7792 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__conb_1_3/HI -0.012f
C7793 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/Q_N -4.33e-20
C7794 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__inv_1_60/Y 0.00442f
C7795 sky130_fd_sc_hd__conb_1_5/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 1.08e-20
C7796 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_31/LO 8.81e-20
C7797 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF18.Q 3.52e-20
C7798 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# 2.84e-32
C7799 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_941_21# -1.62e-20
C7800 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# -2.28e-19
C7801 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 2.21e-19
C7802 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__conb_1_19/HI 6.41e-19
C7803 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 0.00106f
C7804 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_1_48/Y 9.71e-19
C7805 sky130_fd_sc_hd__dfbbn_1_39/a_557_413# V_LOW 3.56e-20
C7806 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_66/A 0.0398f
C7807 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 2.2e-19
C7808 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0963f
C7809 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0076f
C7810 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.043f
C7811 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00496f
C7812 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 0.0218f
C7813 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.0277f
C7814 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_1_29/Y 0.0365f
C7815 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_20/Y 0.0371f
C7816 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 1.44e-20
C7817 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_791_47# 5.45e-20
C7818 sky130_fd_sc_hd__inv_16_41/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 0.331f
C7819 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 3.53e-20
C7820 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.27e-20
C7821 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 1.46e-20
C7822 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__conb_1_33/HI 0.0198f
C7823 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0.00123f
C7824 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_9/Y 0.135f
C7825 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_31/HI 2.22e-20
C7826 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_31/Y 2.25e-20
C7827 sky130_fd_sc_hd__inv_16_51/Y sky130_fd_sc_hd__inv_16_55/Y 0.295f
C7828 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__inv_1_27/Y 1.07e-20
C7829 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 5.16e-19
C7830 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/Q_N 5.16e-19
C7831 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# Reset 0.00104f
C7832 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__conb_1_23/HI 0.00462f
C7833 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# 0.00115f
C7834 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# CLOCK_GEN.SR_Op.Q 5.17e-19
C7835 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.0241f
C7836 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0.00601f
C7837 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 1.23e-20
C7838 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# sky130_fd_sc_hd__conb_1_2/HI 5.88e-20
C7839 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00178f
C7840 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 0.0398f
C7841 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.14f
C7842 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_19/A 0.116f
C7843 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -7.6e-19
C7844 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# -0.00125f
C7845 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -9.88e-20
C7846 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# -0.00228f
C7847 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0236f
C7848 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.00112f
C7849 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0142f
C7850 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__conb_1_25/HI 4.11e-22
C7851 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_1_32/Y 0.0267f
C7852 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__conb_1_11/HI 0.00788f
C7853 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 0.00184f
C7854 sky130_fd_sc_hd__inv_1_22/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 0.107f
C7855 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# -0.00107f
C7856 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# -3.46e-20
C7857 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# 6.21e-21
C7858 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_1_69/Y 7.22e-21
C7859 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# -9.32e-20
C7860 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 3.03e-21
C7861 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 6.89e-19
C7862 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 8.98e-19
C7863 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 0.00829f
C7864 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__inv_1_38/Y 0.00192f
C7865 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_50/Y 2.2e-20
C7866 sky130_fd_sc_hd__conb_1_47/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 1.99e-20
C7867 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_47/a_381_47# 2.34e-20
C7868 sky130_fd_sc_hd__inv_1_43/Y RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0148f
C7869 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_36/Y 0.0407f
C7870 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# V_LOW 0.0438f
C7871 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 0.00367f
C7872 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# -0.00144f
C7873 RISING_COUNTER.COUNT_SUB_DFF0.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.8f
C7874 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 1.97e-21
C7875 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# V_LOW -0.00102f
C7876 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# V_LOW -0.00389f
C7877 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 3.3e-19
C7878 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# -2.57e-20
C7879 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_59/Y 0.0302f
C7880 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# V_LOW 0.0238f
C7881 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# -0.223f
C7882 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__conb_1_46/HI 0.228f
C7883 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# sky130_fd_sc_hd__inv_1_60/Y 0.00185f
C7884 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_28/HI 4.42e-19
C7885 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0246f
C7886 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# Reset 0.048f
C7887 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_1_44/A 0.00347f
C7888 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_381_47# 0.0352f
C7889 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_1_60/Y 2.12e-21
C7890 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# -1.64e-19
C7891 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# V_LOW 0.0139f
C7892 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_1_48/Y 0.0181f
C7893 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00202f
C7894 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 4.78e-19
C7895 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_35/Y 3e-19
C7896 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.00505f
C7897 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.0085f
C7898 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0397f
C7899 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_55/Y 0.00747f
C7900 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nor2_1_0/Y 0.0555f
C7901 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 0.0636f
C7902 sky130_fd_sc_hd__inv_1_30/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00194f
C7903 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 2.85e-20
C7904 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 2.85e-20
C7905 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.027f
C7906 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 6.82e-20
C7907 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 2.52e-19
C7908 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 9.75e-19
C7909 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 1.68e-19
C7910 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_40/Y 0.0308f
C7911 sky130_fd_sc_hd__conb_1_22/HI V_LOW 0.123f
C7912 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0335f
C7913 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__inv_1_43/Y 0.0323f
C7914 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 0.00413f
C7915 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_1_37/Y 8.24e-20
C7916 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_37/HI 0.00698f
C7917 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.03f
C7918 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 1.86e-20
C7919 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# V_LOW 0.0297f
C7920 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 2.22e-20
C7921 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 3.2e-21
C7922 sky130_fd_sc_hd__inv_1_21/Y Reset 0.0165f
C7923 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0121f
C7924 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.15e-19
C7925 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 3.05e-20
C7926 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 7.17e-20
C7927 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0869f
C7928 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.71e-19
C7929 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 0.00181f
C7930 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 4.63e-19
C7931 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 2.02e-19
C7932 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_51/Y 0.184f
C7933 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0874f
C7934 sky130_fd_sc_hd__inv_1_10/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 1.17e-20
C7935 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__conb_1_25/HI 0.00112f
C7936 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__inv_1_28/Y 0.00117f
C7937 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# V_LOW 4.8e-20
C7938 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__conb_1_6/HI 5.52e-19
C7939 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_16_41/Y 0.196f
C7940 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# 6.75e-19
C7941 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# V_LOW 0.0147f
C7942 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_557_413# 4.16e-19
C7943 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_65/Y 0.0109f
C7944 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/Q_N -4.24e-20
C7945 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 7.01e-19
C7946 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_791_47# 7.04e-19
C7947 sky130_fd_sc_hd__inv_1_46/A FULL_COUNTER.COUNT_SUB_DFF0.Q 8.32e-19
C7948 sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_15/A 0.168f
C7949 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 1.76e-19
C7950 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# sky130_fd_sc_hd__inv_1_38/Y 6.84e-22
C7951 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__inv_1_36/Y 1.01e-20
C7952 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_1/Y 0.024f
C7953 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 0.00407f
C7954 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# -0.0047f
C7955 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# -0.00125f
C7956 sky130_fd_sc_hd__inv_16_48/Y CLOCK_GEN.SR_Op.Q 0.023f
C7957 sky130_fd_sc_hd__conb_1_7/HI V_LOW 0.315f
C7958 FULL_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 1.36f
C7959 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__conb_1_44/LO 3.58e-20
C7960 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# sky130_fd_sc_hd__inv_16_41/Y 4.63e-20
C7961 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00597f
C7962 sky130_fd_sc_hd__inv_16_40/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0196f
C7963 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# V_LOW 2.94e-20
C7964 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 1.05e-19
C7965 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 2.6e-20
C7966 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# -0.00141f
C7967 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_16_40/Y 0.00641f
C7968 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.4e-21
C7969 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_24/Y 7.14e-20
C7970 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_35/Y 0.0954f
C7971 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 1.54e-20
C7972 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00152f
C7973 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 2.43e-20
C7974 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00389f
C7975 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__inv_1_59/Y 0.00713f
C7976 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# V_LOW 0.00946f
C7977 sky130_fd_sc_hd__conb_1_46/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.95e-20
C7978 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.1e-20
C7979 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_45/LO 0.00103f
C7980 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# -2.52e-19
C7981 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -0.0116f
C7982 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 2.84e-32
C7983 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 0.732f
C7984 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_16/HI 0.103f
C7985 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0232f
C7986 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__conb_1_17/HI 9.28e-22
C7987 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_23/HI 0.113f
C7988 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# Reset 0.00291f
C7989 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# sky130_fd_sc_hd__inv_1_44/A 4.96e-19
C7990 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# V_LOW 1.79e-20
C7991 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_1_7/Y 1.57e-20
C7992 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# V_LOW 3.56e-20
C7993 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.51e-19
C7994 sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.00731f
C7995 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__inv_1_34/Y 9.59e-20
C7996 sky130_fd_sc_hd__conb_1_41/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00163f
C7997 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# -6.23e-21
C7998 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# -6.22e-19
C7999 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_381_47# -4.37e-20
C8000 sky130_fd_sc_hd__dfbbn_1_44/Q_N RISING_COUNTER.COUNT_SUB_DFF4.Q 1.04e-19
C8001 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 2.01e-20
C8002 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 4.71e-20
C8003 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.1e-21
C8004 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_1_63/Y 5.2e-20
C8005 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 9.37e-20
C8006 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.02e-21
C8007 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 0.00115f
C8008 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_1_46/A 0.0717f
C8009 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__inv_1_37/Y 1.17e-19
C8010 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.71e-19
C8011 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# -0.0309f
C8012 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_557_413# -3.67e-20
C8013 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__inv_1_27/Y 5.85e-22
C8014 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__inv_1_24/A 1.61e-19
C8015 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# V_LOW 0.0126f
C8016 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__inv_1_38/Y 0.00116f
C8017 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI 7.33e-19
C8018 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 0.00127f
C8019 sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF6.Q 0.434f
C8020 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_56/Y 0.0423f
C8021 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_46/A 7.6e-21
C8022 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.46e-19
C8023 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.254f
C8024 sky130_fd_sc_hd__nand2_8_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.8e-20
C8025 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# V_LOW 0.00734f
C8026 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0274f
C8027 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.51e-19
C8028 RISING_COUNTER.COUNT_SUB_DFF1.Q V_HIGH 1.43f
C8029 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/Q_N -4.24e-20
C8030 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/Q_N -9.56e-20
C8031 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_8_0/A 1.35e-19
C8032 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00551f
C8033 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_42/LO 0.0141f
C8034 sky130_fd_sc_hd__conb_1_22/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 7.81e-20
C8035 sky130_fd_sc_hd__inv_1_32/Y FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00397f
C8036 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_9/A 4.53e-19
C8037 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.09e-19
C8038 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 0.00114f
C8039 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# 5.39e-19
C8040 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# V_LOW 2.94e-20
C8041 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 2.79e-20
C8042 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# -0.00146f
C8043 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# -3.65e-19
C8044 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_1_42/Y 4.44e-20
C8045 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# V_LOW -0.00446f
C8046 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0143f
C8047 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.32e-20
C8048 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0379f
C8049 sky130_fd_sc_hd__conb_1_44/HI V_LOW 0.123f
C8050 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0089f
C8051 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0124f
C8052 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# 0.00387f
C8053 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_381_47# -2.53e-20
C8054 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_66/A 0.00144f
C8055 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_33/Y 0.202f
C8056 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_46/A 0.0444f
C8057 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/Q_N 0.00266f
C8058 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_17/HI 6.4e-19
C8059 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_22/A 0.00528f
C8060 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.67e-21
C8061 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# 5.26e-22
C8062 sky130_fd_sc_hd__dfbbn_1_11/Q_N V_LOW -2.68e-19
C8063 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 5.73e-20
C8064 Reset sky130_fd_sc_hd__conb_1_37/HI 0.215f
C8065 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__conb_1_37/HI 0.0147f
C8066 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00392f
C8067 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# V_LOW -0.00266f
C8068 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_51/Y 0.0895f
C8069 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 9.04e-20
C8070 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# -1.76e-19
C8071 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__inv_1_41/Y 0.00468f
C8072 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__conb_1_5/HI 3.91e-20
C8073 sky130_fd_sc_hd__conb_1_51/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 4.75e-19
C8074 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 3.77e-20
C8075 sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16_50/A 0.00271f
C8076 sky130_fd_sc_hd__inv_16_51/A sky130_fd_sc_hd__inv_16_48/A 0.56f
C8077 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_44/A 0.0406f
C8078 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_23/HI 0.0238f
C8079 sky130_fd_sc_hd__inv_16_24/Y V_LOW 0.0903f
C8080 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_8/Y 0.00772f
C8081 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_44/HI 6.85e-20
C8082 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 1.8e-21
C8083 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 3.77e-20
C8084 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_17/HI -5.71e-19
C8085 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_18/A 5.2e-20
C8086 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# sky130_fd_sc_hd__conb_1_34/HI 0.0017f
C8087 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0541f
C8088 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__conb_1_20/HI 5.58e-21
C8089 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0314f
C8090 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 1.48e-19
C8091 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.0613f
C8092 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_647_21# -8.61e-20
C8093 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# -1.63e-19
C8094 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_19/HI -0.00469f
C8095 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__conb_1_30/HI -2.07e-19
C8096 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 0.00322f
C8097 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00322f
C8098 sky130_fd_sc_hd__nand3_1_1/a_193_47# sky130_fd_sc_hd__inv_1_64/Y 7.46e-19
C8099 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_21/Y 2.81e-19
C8100 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 1.23e-21
C8101 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_50/HI 0.472f
C8102 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_67/A 0.0364f
C8103 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0215f
C8104 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00356f
C8105 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__conb_1_21/HI -0.00581f
C8106 sky130_fd_sc_hd__conb_1_5/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 1.53e-19
C8107 sky130_fd_sc_hd__conb_1_29/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0127f
C8108 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0014f
C8109 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0044f
C8110 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_31/Y 0.00172f
C8111 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.61e-19
C8112 sky130_fd_sc_hd__nand2_8_7/a_27_47# Reset 0.00244f
C8113 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_2_0/A 1.65e-19
C8114 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_24/HI 0.0152f
C8115 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 0.0754f
C8116 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__inv_1_38/Y 0.21f
C8117 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_19/A 0.0126f
C8118 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_7/Y 0.26f
C8119 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_51/A 0.00238f
C8120 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00215f
C8121 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/Q_N 4.28e-20
C8122 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__conb_1_16/HI 6e-19
C8123 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_1_22/Y 7.13e-19
C8124 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__inv_1_62/Y 0.0154f
C8125 sky130_fd_sc_hd__inv_16_29/Y sky130_fd_sc_hd__inv_16_28/Y 0.0113f
C8126 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 4.6e-20
C8127 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 1.3e-19
C8128 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 3.03e-21
C8129 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 8.98e-19
C8130 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 6.89e-19
C8131 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# -1.65e-19
C8132 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# -5.16e-20
C8133 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 7.3e-19
C8134 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_24/A 0.378f
C8135 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.01e-20
C8136 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0416f
C8137 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0137f
C8138 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__inv_1_36/Y 6.66e-20
C8139 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/Q_N -9.56e-20
C8140 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_25/HI 0.035f
C8141 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# -1.44e-20
C8142 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0253f
C8143 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 5.8e-20
C8144 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00147f
C8145 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 3.4e-20
C8146 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# V_LOW 1.38e-19
C8147 FULL_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0255f
C8148 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# -0.00393f
C8149 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_557_413# -0.0012f
C8150 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__conb_1_4/HI 0.0215f
C8151 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 8.59e-20
C8152 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__inv_16_42/Y 0.00289f
C8153 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.0243f
C8154 sky130_fd_sc_hd__conb_1_17/HI V_LOW 0.219f
C8155 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_26/Y 6.69e-21
C8156 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_51/A 0.00774f
C8157 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.12e-19
C8158 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_47/Y 0.152f
C8159 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_473_413# -0.00985f
C8160 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_647_21# -6.43e-20
C8161 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__conb_1_23/HI 0.00482f
C8162 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_557_413# -0.0012f
C8163 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# -0.0256f
C8164 sky130_fd_sc_hd__inv_1_62/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0886f
C8165 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 3.56e-19
C8166 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__inv_1_61/Y 0.00207f
C8167 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# V_LOW 0.00883f
C8168 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 2.2e-20
C8169 sky130_fd_sc_hd__inv_16_6/A Reset 0.318f
C8170 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__nand2_8_4/Y 6.56e-20
C8171 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/Q_N -9.56e-20
C8172 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__conb_1_17/HI -3.23e-20
C8173 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.03e-21
C8174 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.3e-19
C8175 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0.0112f
C8176 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0.00104f
C8177 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 0.00215f
C8178 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_1_25/Y 3.69e-19
C8179 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 2.62e-20
C8180 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# V_LOW 0.00245f
C8181 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 0.0514f
C8182 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16_52/A 0.208f
C8183 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_581_47# -7.91e-19
C8184 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# -0.0567f
C8185 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 3.43e-19
C8186 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# -0.00336f
C8187 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# -3.79e-20
C8188 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.117f
C8189 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.0349f
C8190 sky130_fd_sc_hd__conb_1_25/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 5e-20
C8191 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__conb_1_19/HI 0.00689f
C8192 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 4.12e-20
C8193 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 4.12e-20
C8194 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.006f
C8195 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.0108f
C8196 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# 8.69e-19
C8197 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 2.54e-19
C8198 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.38e-19
C8199 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_8_9/A 0.0757f
C8200 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -3.48e-20
C8201 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 0.0172f
C8202 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# V_LOW 0.0249f
C8203 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 7.69e-20
C8204 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__conb_1_21/HI 5.27e-20
C8205 sky130_fd_sc_hd__dfbbn_1_47/Q_N V_LOW -2.68e-19
C8206 sky130_fd_sc_hd__conb_1_13/LO V_LOW 0.0859f
C8207 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__inv_1_31/Y 0.00146f
C8208 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.13e-19
C8209 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 0.00553f
C8210 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 0.0306f
C8211 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__conb_1_37/HI 0.236f
C8212 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand3_1_1/Y 0.00205f
C8213 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_1_37/Y 4.43e-21
C8214 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# Reset 0.0252f
C8215 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00158f
C8216 sky130_fd_sc_hd__inv_1_42/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 3.8e-19
C8217 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# V_LOW 1.38e-19
C8218 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_10/HI 0.0181f
C8219 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__nand2_8_9/A 6.86e-21
C8220 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 7.01e-19
C8221 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_791_47# 7.04e-19
C8222 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 9.05e-19
C8223 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.003f
C8224 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 8.4e-21
C8225 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 6.66e-19
C8226 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_29/HI -0.00108f
C8227 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00995f
C8228 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00119f
C8229 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.00575f
C8230 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 4.27e-20
C8231 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__conb_1_25/HI 0.0138f
C8232 sky130_fd_sc_hd__inv_1_67/Y Reset 0.0176f
C8233 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.41e-19
C8234 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 1.02e-19
C8235 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_43/HI 0.00793f
C8236 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# -3.86e-20
C8237 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_941_21# -8.98e-20
C8238 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# Reset 0.0155f
C8239 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.166f
C8240 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_25/LO 2.62e-19
C8241 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 2.52e-21
C8242 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.65e-19
C8243 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# -6.43e-20
C8244 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# -5.78e-20
C8245 sky130_fd_sc_hd__inv_1_53/Y V_LOW 0.0567f
C8246 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# sky130_fd_sc_hd__conb_1_4/HI -0.0119f
C8247 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__conb_1_37/HI -6.23e-19
C8248 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.96e-19
C8249 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 1.86e-21
C8250 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 3.37e-20
C8251 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 0.00347f
C8252 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_44/A 0.00398f
C8253 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00109f
C8254 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.00479f
C8255 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 9.28e-19
C8256 V_SENSE CLOCK_GEN.SR_Op.Q 1.19f
C8257 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# -1.69e-19
C8258 sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.106f
C8259 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -5.42e-19
C8260 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# 5.32e-19
C8261 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 4.56e-21
C8262 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 1.65e-19
C8263 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 2.69e-20
C8264 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# V_LOW 1.79e-20
C8265 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 1.07e-20
C8266 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0354f
C8267 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 0.0922f
C8268 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.01e-21
C8269 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__conb_1_46/HI 1.36e-20
C8270 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 1.07e-19
C8271 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# V_LOW 0.0191f
C8272 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_23/Y 6.96e-19
C8273 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__conb_1_18/HI 0.0121f
C8274 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_44/A 8.51e-20
C8275 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_28/HI 0.255f
C8276 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 0.0331f
C8277 FULL_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 0.325f
C8278 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_473_413# 1.62e-19
C8279 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__conb_1_26/HI 0.038f
C8280 sky130_fd_sc_hd__inv_16_40/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.045f
C8281 sky130_fd_sc_hd__inv_16_41/Y CLOCK_GEN.SR_Op.Q 4.08e-20
C8282 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# -0.00512f
C8283 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# -0.00117f
C8284 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 4.57e-20
C8285 sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__inv_1_19/Y 0.03f
C8286 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_17/HI 0.15f
C8287 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__conb_1_19/HI -2.17e-19
C8288 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0148f
C8289 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__conb_1_11/HI -0.00643f
C8290 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0335f
C8291 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.109f
C8292 V_SENSE sky130_fd_sc_hd__inv_1_63/Y 7.8e-19
C8293 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__inv_1_26/Y 0.00808f
C8294 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# V_LOW -0.00336f
C8295 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# 8.32e-19
C8296 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# V_LOW 0.01f
C8297 sky130_fd_sc_hd__dfbbn_1_15/Q_N FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0277f
C8298 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_24/LO 3.72e-20
C8299 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__conb_1_21/HI -2.17e-19
C8300 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 0.111f
C8301 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 1.82e-19
C8302 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 2.87e-20
C8303 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_3/HI 0.0249f
C8304 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00138f
C8305 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_6/HI 0.2f
C8306 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 2.32e-19
C8307 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0273f
C8308 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0569f
C8309 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_1_37/Y 1.42e-19
C8310 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# 3.38e-20
C8311 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_51/Y 1.46e-21
C8312 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 1.47e-19
C8313 sky130_fd_sc_hd__dfbbn_1_44/Q_N FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00841f
C8314 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# Reset 0.00539f
C8315 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_891_329# -3.85e-20
C8316 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# -3.48e-20
C8317 sky130_fd_sc_hd__inv_1_4/Y V_LOW 0.136f
C8318 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__conb_1_26/LO 3.22e-20
C8319 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__conb_1_10/HI 0.00248f
C8320 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_65/A 1.6e-19
C8321 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.37e-20
C8322 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 5.28e-19
C8323 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 2.39e-20
C8324 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.18e-20
C8325 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_24/LO 4.69e-21
C8326 sky130_fd_sc_hd__conb_1_45/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 8.81e-21
C8327 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00606f
C8328 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_26/HI 1.65e-20
C8329 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0167f
C8330 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_32/Y 6.74e-22
C8331 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__inv_1_62/Y 1.21e-20
C8332 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__inv_1_50/Y 0.00506f
C8333 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_50/HI 0.108f
C8334 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# -8.61e-20
C8335 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_29/A 1.03e-19
C8336 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_44/A 0.00117f
C8337 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# sky130_fd_sc_hd__conb_1_44/HI 0.0049f
C8338 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# sky130_fd_sc_hd__conb_1_43/HI 6.58e-19
C8339 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.33e-19
C8340 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0.0138f
C8341 sky130_fd_sc_hd__inv_1_39/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.04e-22
C8342 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# -1.06e-19
C8343 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00236f
C8344 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# Reset 3.02e-19
C8345 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0216f
C8346 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_55/Y 0.228f
C8347 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.18e-19
C8348 sky130_fd_sc_hd__fill_8_858/VPB V_LOW 0.797f
C8349 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# CLOCK_GEN.SR_Op.Q 1.71e-19
C8350 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00143f
C8351 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 1.67e-19
C8352 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# sky130_fd_sc_hd__conb_1_37/HI -0.00265f
C8353 sky130_fd_sc_hd__nand2_8_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 8.11e-21
C8354 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.12f
C8355 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 3.77e-19
C8356 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 4.04e-19
C8357 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_581_47# -7.91e-19
C8358 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_1_22/Y 0.0026f
C8359 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.83e-20
C8360 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 3.01e-20
C8361 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# 2.1e-20
C8362 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 6.24e-21
C8363 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_6/HI 1.58e-20
C8364 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_30/Y 0.0465f
C8365 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 0.0015f
C8366 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 6.58e-20
C8367 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0228f
C8368 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q -2.49e-20
C8369 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 1.65e-21
C8370 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.05f
C8371 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# 1.19e-19
C8372 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__inv_1_36/Y 0.00464f
C8373 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 5.4e-19
C8374 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.78e-21
C8375 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# -0.00834f
C8376 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# -5.02e-19
C8377 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_24/A 0.00284f
C8378 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_16/HI 0.00408f
C8379 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_1_25/Y 1.89e-21
C8380 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0411f
C8381 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 8.79e-22
C8382 sky130_fd_sc_hd__inv_1_9/Y V_LOW 0.369f
C8383 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 2.76e-20
C8384 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# -4.66e-20
C8385 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# -3.79e-20
C8386 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# V_LOW 3.56e-20
C8387 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# 0.00307f
C8388 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# V_LOW 0.00508f
C8389 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_16/HI 0.112f
C8390 sky130_fd_sc_hd__dfbbn_1_20/a_581_47# sky130_fd_sc_hd__conb_1_18/HI 3.73e-19
C8391 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# V_LOW 1.69e-19
C8392 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0249f
C8393 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__conb_1_30/HI 0.0116f
C8394 sky130_fd_sc_hd__conb_1_9/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 7.35e-20
C8395 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_40/Y 3.55e-21
C8396 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 3.83e-19
C8397 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# 0.0018f
C8398 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 1.9e-19
C8399 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# sky130_fd_sc_hd__inv_1_12/Y 1.5e-21
C8400 sky130_fd_sc_hd__conb_1_39/LO Reset 1.54e-19
C8401 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__nand2_8_4/Y 4.53e-21
C8402 sky130_fd_sc_hd__inv_1_57/Y V_LOW 0.189f
C8403 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_647_21# -0.00499f
C8404 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 3.45e-19
C8405 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_16_2/Y 1.51e-20
C8406 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0104f
C8407 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.0439f
C8408 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# V_LOW -2.48e-19
C8409 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# sky130_fd_sc_hd__conb_1_11/HI 1.1e-19
C8410 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0354f
C8411 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0234f
C8412 sky130_fd_sc_hd__inv_16_15/Y sky130_fd_sc_hd__inv_16_15/A 0.15f
C8413 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# V_LOW -1.39e-35
C8414 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00146f
C8415 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_44/A 6.48e-19
C8416 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__conb_1_18/LO 0.00434f
C8417 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 8.92e-19
C8418 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_67/A 3.93e-21
C8419 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 9.26e-20
C8420 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_2_0/A 0.125f
C8421 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0136f
C8422 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_1_44/A 0.0162f
C8423 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.18e-20
C8424 sky130_fd_sc_hd__inv_1_19/A V_LOW 0.973f
C8425 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 1.55e-21
C8426 sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__inv_1_56/A 5.96e-19
C8427 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.33e-19
C8428 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# -3.46e-20
C8429 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# V_LOW 1.38e-19
C8430 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__conb_1_12/HI 3.01e-21
C8431 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 6.21e-20
C8432 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 2.93e-20
C8433 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 3.94e-19
C8434 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# -0.00183f
C8435 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.39e-19
C8436 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_25/HI 3.41e-19
C8437 sky130_fd_sc_hd__conb_1_33/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 2.55e-19
C8438 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 1.43e-19
C8439 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 1.91e-20
C8440 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0197f
C8441 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__conb_1_50/HI 4.09e-19
C8442 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_581_47# -7.91e-19
C8443 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00249f
C8444 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.22e-19
C8445 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_67/A 0.129f
C8446 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# V_LOW 0.0057f
C8447 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 0.00152f
C8448 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.16e-19
C8449 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# V_LOW -0.00483f
C8450 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# CLOCK_GEN.SR_Op.Q 8.81e-19
C8451 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 2.4e-20
C8452 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 0.00453f
C8453 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 4.95e-19
C8454 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 0.0109f
C8455 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 5.15e-19
C8456 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_64/Y 0.003f
C8457 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0138f
C8458 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0471f
C8459 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 8.66e-21
C8460 sky130_fd_sc_hd__conb_1_29/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0205f
C8461 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 2.66e-19
C8462 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00708f
C8463 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# 5.54e-20
C8464 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# 5.86e-21
C8465 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.53e-21
C8466 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_581_47# 2.47e-19
C8467 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00709f
C8468 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_9/HI 4.58e-19
C8469 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 2.47e-20
C8470 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# V_LOW 0.0236f
C8471 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_49/Y 0.696f
C8472 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__conb_1_33/HI 1.12e-19
C8473 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_557_413# 8.26e-19
C8474 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 0.0362f
C8475 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.79e-19
C8476 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 6.84e-20
C8477 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.307f
C8478 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# -2.57e-20
C8479 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_1_46/A 9.08e-20
C8480 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# -2.48e-19
C8481 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -0.00151f
C8482 sky130_fd_sc_hd__dfbbn_1_23/Q_N FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0231f
C8483 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__conb_1_31/HI -0.00181f
C8484 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__conb_1_16/HI 0.0155f
C8485 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 8.4e-20
C8486 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -3.24e-20
C8487 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_38/LO 7.4e-19
C8488 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.046f
C8489 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_47/Y 0.142f
C8490 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_19/Y 0.114f
C8491 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_67/A 1.6e-21
C8492 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_891_329# -2.2e-20
C8493 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# -4.1e-19
C8494 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 2.2e-20
C8495 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 0.00335f
C8496 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0387f
C8497 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# V_LOW 0.0137f
C8498 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 0.00125f
C8499 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_33/LO 8.84e-20
C8500 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.0281f
C8501 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 7.85e-20
C8502 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__nand2_8_8/A 2.7e-19
C8503 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_28/HI -0.00114f
C8504 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_581_47# -2.6e-20
C8505 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__nand2_1_2/A 9.87e-21
C8506 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 0.0692f
C8507 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_25/Y 1.15e-19
C8508 sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__conb_1_11/HI 4.43e-20
C8509 sky130_fd_sc_hd__conb_1_26/LO FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.036f
C8510 FULL_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.021f
C8511 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_47/A 0.0134f
C8512 sky130_fd_sc_hd__dfbbn_1_18/Q_N V_LOW -0.00993f
C8513 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__inv_1_49/Y 1.07e-20
C8514 sky130_fd_sc_hd__dfbbn_1_46/Q_N FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0054f
C8515 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_15/Y 2.71e-19
C8516 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 9.28e-19
C8517 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.15e-19
C8518 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 6.4e-19
C8519 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00596f
C8520 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.94e-20
C8521 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_33/Y 1.6e-19
C8522 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0105f
C8523 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__conb_1_20/HI 0.00303f
C8524 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__inv_1_2/Y 9.28e-21
C8525 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.82e-20
C8526 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__inv_1_44/A 1.9e-19
C8527 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1_41/Y 2.43e-19
C8528 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 1.27e-20
C8529 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 2.55e-21
C8530 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_42/Y 0.0402f
C8531 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 7.31e-19
C8532 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__conb_1_25/HI 3.29e-20
C8533 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.0435f
C8534 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# sky130_fd_sc_hd__inv_1_13/Y 9.11e-20
C8535 sky130_fd_sc_hd__inv_1_49/Y V_LOW 0.0218f
C8536 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 4.18e-19
C8537 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__conb_1_0/HI -9.62e-19
C8538 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__conb_1_21/HI 0.00167f
C8539 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__inv_1_12/Y 6.7e-19
C8540 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# V_LOW 3.56e-20
C8541 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 0.347f
C8542 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.71e-19
C8543 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.102f
C8544 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__inv_1_45/Y 0.0108f
C8545 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/Q_N 8.37e-19
C8546 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 6.26e-20
C8547 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.004f
C8548 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_38/Y 0.125f
C8549 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/Q_N 4.46e-21
C8550 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 2.27e-19
C8551 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.95e-19
C8552 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00289f
C8553 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/Q_N 1.15e-19
C8554 FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF7.Q 2.63f
C8555 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 6.86e-19
C8556 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_4/HI 0.00143f
C8557 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__conb_1_6/HI 1.62e-19
C8558 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# V_LOW 0.0144f
C8559 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# -0.0395f
C8560 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# V_LOW 2.94e-20
C8561 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_473_413# 0.0484f
C8562 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__conb_1_33/HI -0.00746f
C8563 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00114f
C8564 sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00101f
C8565 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00236f
C8566 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# -7.17e-20
C8567 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# -1.76e-19
C8568 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# sky130_fd_sc_hd__inv_1_69/Y 3.75e-21
C8569 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0116f
C8570 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_11/LO 0.00206f
C8571 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 8.34e-19
C8572 sky130_fd_sc_hd__conb_1_31/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0141f
C8573 sky130_fd_sc_hd__conb_1_26/HI sky130_fd_sc_hd__conb_1_23/HI 0.0263f
C8574 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_29/HI 1.49e-21
C8575 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00431f
C8576 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_15/HI 0.00463f
C8577 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# -0.00385f
C8578 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 1.38e-20
C8579 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_18/A 0.0277f
C8580 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.05e-19
C8581 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.26e-22
C8582 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# -2.01e-20
C8583 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_6/A 0.0932f
C8584 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 0.00428f
C8585 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_1_36/Y 0.00254f
C8586 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_28/HI -2.07e-19
C8587 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 2.2e-20
C8588 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_20/Y 0.00272f
C8589 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0144f
C8590 sky130_fd_sc_hd__dfbbn_1_35/Q_N V_LOW -0.00509f
C8591 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00149f
C8592 sky130_fd_sc_hd__dfbbn_1_43/Q_N FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.025f
C8593 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 8.16e-19
C8594 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_19/LO 1.95e-20
C8595 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.08e-19
C8596 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__conb_1_2/HI 1.98e-19
C8597 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00115f
C8598 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 9.94e-20
C8599 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# sky130_fd_sc_hd__inv_1_33/Y 0.00164f
C8600 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 0.00363f
C8601 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# V_LOW 0.0112f
C8602 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__conb_1_19/HI 3.01e-21
C8603 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# Reset 0.0387f
C8604 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__conb_1_23/HI 5.57e-21
C8605 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 4.15e-22
C8606 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_891_329# -0.00159f
C8607 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# -0.00942f
C8608 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_20/Y 0.0171f
C8609 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# 1.89e-19
C8610 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0024f
C8611 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# -0.00869f
C8612 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 2.64e-19
C8613 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/Q_N -4.33e-20
C8614 sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF15.Q 0.133f
C8615 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__conb_1_30/HI 9.42e-19
C8616 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_60/Y 0.185f
C8617 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.013f
C8618 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 9.27e-19
C8619 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__inv_1_9/Y 1.98e-20
C8620 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_67/A 1.85e-20
C8621 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_14/Y -0.00363f
C8622 FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 0.497f
C8623 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.0114f
C8624 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 5.4e-20
C8625 sky130_fd_sc_hd__inv_16_40/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0335f
C8626 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_26/Y 0.00173f
C8627 sky130_fd_sc_hd__dfbbn_1_18/Q_N RISING_COUNTER.COUNT_SUB_DFF13.Q 1.56e-20
C8628 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_46/A 2.26e-21
C8629 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.85e-20
C8630 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0051f
C8631 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# sky130_fd_sc_hd__conb_1_11/HI 1.1e-21
C8632 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 1.76e-20
C8633 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 3.48e-19
C8634 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 6.77e-20
C8635 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 1.14e-19
C8636 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.92e-20
C8637 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.34e-19
C8638 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00616f
C8639 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_29/HI 0.00271f
C8640 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__conb_1_50/HI 4.24e-19
C8641 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__nand2_8_8/A 7.18e-19
C8642 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# sky130_fd_sc_hd__conb_1_6/HI 0.00183f
C8643 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1_44/LO 0.00126f
C8644 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# V_LOW 0.01f
C8645 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.00776f
C8646 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/a_193_47# 5.58e-20
C8647 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0.00138f
C8648 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 0.0122f
C8649 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.94e-20
C8650 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__inv_1_28/Y 0.00506f
C8651 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_29/Y 0.0964f
C8652 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_2_0/A 0.0616f
C8653 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_1_21/Y 0.00179f
C8654 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/Q_N -6.48e-19
C8655 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_5/A 0.00643f
C8656 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# -0.02f
C8657 sky130_fd_sc_hd__nand3_1_0/Y V_LOW 1.63f
C8658 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0265f
C8659 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00213f
C8660 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00238f
C8661 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 1.38e-20
C8662 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 2.26e-19
C8663 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 6.57e-19
C8664 sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0501f
C8665 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.7e-20
C8666 sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__inv_1_50/Y 0.00148f
C8667 sky130_fd_sc_hd__inv_1_41/Y V_LOW 0.281f
C8668 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 2.75e-19
C8669 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__conb_1_23/LO 9.95e-20
C8670 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 1.47e-20
C8671 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 3.71e-19
C8672 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__conb_1_2/HI 1.51e-19
C8673 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# V_LOW 5.79e-19
C8674 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/Q_N 5.21e-19
C8675 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_1_33/Y 0.00345f
C8676 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_1_5/Y 0.0888f
C8677 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 2e-20
C8678 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__inv_16_42/Y 1.18e-19
C8679 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 2.51e-20
C8680 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 5.3e-22
C8681 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 1.91e-20
C8682 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 1.25e-19
C8683 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# Reset 0.0624f
C8684 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.79e-20
C8685 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# CLOCK_GEN.SR_Op.Q 0.287f
C8686 sky130_fd_sc_hd__conb_1_51/HI V_LOW 0.0993f
C8687 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# V_LOW 0.0264f
C8688 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__conb_1_23/HI -6.57e-19
C8689 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.99e-20
C8690 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__inv_1_1/Y 7.97e-21
C8691 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# -0.00552f
C8692 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0158f
C8693 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.262f
C8694 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0827f
C8695 sky130_fd_sc_hd__dfbbn_1_12/a_581_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 3.35e-19
C8696 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# -0.00107f
C8697 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# -2.53e-20
C8698 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00782f
C8699 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0366f
C8700 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 3.71e-20
C8701 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# V_LOW 1.45e-19
C8702 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 0.00223f
C8703 sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__inv_1_47/Y 0.00878f
C8704 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_65/A 1.82e-19
C8705 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_24/Y 2.55e-19
C8706 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.0666f
C8707 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.0398f
C8708 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0453f
C8709 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# 0.00167f
C8710 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_8/Y 0.00535f
C8711 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__inv_16_41/Y 0.00112f
C8712 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_61/Y 0.187f
C8713 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_47/Y 6.96e-19
C8714 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__conb_1_4/HI 2.52e-19
C8715 sky130_fd_sc_hd__conb_1_12/LO V_LOW 0.0952f
C8716 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_16_29/Y 0.00427f
C8717 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 3.41e-19
C8718 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# 1.69e-20
C8719 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_1_38/Y 0.00331f
C8720 FULL_COUNTER.COUNT_SUB_DFF19.Q V_LOW 4.67f
C8721 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 1e-20
C8722 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__inv_1_69/Y 0.0011f
C8723 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00769f
C8724 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__conb_1_26/HI 0.043f
C8725 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# -6.23e-21
C8726 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# -0.00502f
C8727 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__conb_1_47/HI 1.36e-19
C8728 RISING_COUNTER.COUNT_SUB_DFF7.Q V_LOW 2.27f
C8729 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_49/Y 5.97e-20
C8730 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__inv_2_0/A 0.0185f
C8731 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 3.83e-19
C8732 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 3.4e-20
C8733 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_19/Y 0.114f
C8734 sky130_fd_sc_hd__conb_1_33/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00101f
C8735 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16_51/Y 0.191f
C8736 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_44/A 0.0018f
C8737 sky130_fd_sc_hd__fill_8_927/VPB V_LOW 0.797f
C8738 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 1.76e-19
C8739 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_23/HI 0.147f
C8740 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/Q_N -4.78e-20
C8741 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_8_0/A 1.11e-19
C8742 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__conb_1_15/HI 0.0116f
C8743 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__conb_1_48/LO 9.76e-21
C8744 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 4.13e-19
C8745 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0301f
C8746 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/Q_N 2.3e-21
C8747 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -0.00953f
C8748 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_891_329# -2.2e-20
C8749 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 1.25e-19
C8750 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_1/LO 0.00813f
C8751 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 7.63e-20
C8752 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 1.28e-19
C8753 sky130_fd_sc_hd__fill_8_854/VPB V_LOW 0.797f
C8754 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__conb_1_15/HI 0.0083f
C8755 sky130_fd_sc_hd__conb_1_29/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0128f
C8756 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 6.18e-19
C8757 sky130_fd_sc_hd__inv_16_6/A FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0299f
C8758 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0411f
C8759 sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF7.Q 0.109f
C8760 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# -0.14f
C8761 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1_25/HI 0.0399f
C8762 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# V_LOW -0.00389f
C8763 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__conb_1_39/HI 8.3e-20
C8764 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# CLOCK_GEN.SR_Op.Q 0.00252f
C8765 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# -0.00144f
C8766 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# V_LOW 0.00665f
C8767 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_20/Y 0.01f
C8768 sky130_fd_sc_hd__conb_1_10/HI V_LOW 0.0254f
C8769 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0449f
C8770 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# V_LOW 0.0108f
C8771 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# V_LOW -0.00389f
C8772 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_1_40/Y 9.93e-21
C8773 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_1_25/Y 1.46e-20
C8774 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.12f
C8775 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_60/Y 6.52e-21
C8776 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.018f
C8777 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_7/HI 0.0187f
C8778 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# -0.00141f
C8779 sky130_fd_sc_hd__dfbbn_1_25/Q_N FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00208f
C8780 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0384f
C8781 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0314f
C8782 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# V_LOW -1.53e-19
C8783 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__conb_1_37/HI 1.31e-20
C8784 sky130_fd_sc_hd__inv_1_5/Y V_LOW 0.388f
C8785 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.49e-21
C8786 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# V_LOW -9.15e-19
C8787 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# sky130_fd_sc_hd__inv_1_39/Y 2.62e-19
C8788 sky130_fd_sc_hd__inv_1_24/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 1.58e-20
C8789 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.45e-19
C8790 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_64/A 0.866f
C8791 sky130_fd_sc_hd__inv_16_6/A FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.109f
C8792 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 2.16e-19
C8793 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# sky130_fd_sc_hd__inv_16_40/Y 0.00472f
C8794 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 1.41f
C8795 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 0.0226f
C8796 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_39/Y 0.0375f
C8797 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/Q_N 1.18e-19
C8798 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 0.00302f
C8799 sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__inv_16_40/Y 0.145f
C8800 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 2.62e-19
C8801 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_1_46/A 0.00452f
C8802 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__inv_1_69/Y 4.54e-19
C8803 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# sky130_fd_sc_hd__conb_1_26/HI 4.8e-19
C8804 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 8.71e-21
C8805 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# V_LOW -0.0266f
C8806 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.25e-21
C8807 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_45/Y 7.86e-21
C8808 sky130_fd_sc_hd__inv_1_29/Y V_LOW 0.0552f
C8809 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# sky130_fd_sc_hd__conb_1_47/HI -2.6e-20
C8810 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 6.53e-20
C8811 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_28/Y 9.49e-19
C8812 sky130_fd_sc_hd__conb_1_13/HI FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0226f
C8813 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# 9.67e-20
C8814 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_891_329# -2.2e-20
C8815 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# -4.1e-19
C8816 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0841f
C8817 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__conb_1_17/LO 0.0689f
C8818 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_16_2/Y 0.299f
C8819 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_1_44/A 4.56e-19
C8820 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 3.54e-20
C8821 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0644f
C8822 sky130_fd_sc_hd__conb_1_2/LO FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00204f
C8823 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# V_LOW -0.00266f
C8824 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 0.0199f
C8825 V_SENSE sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 7.27e-20
C8826 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 7.39e-20
C8827 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 8.97e-20
C8828 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 7.39e-20
C8829 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.0127f
C8830 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 8.97e-20
C8831 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# -0.00592f
C8832 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# 1.42e-32
C8833 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_16_19/Y 9.23e-19
C8834 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_2_0/A 3.38e-19
C8835 V_SENSE sky130_fd_sc_hd__inv_16_8/A 0.285f
C8836 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0377f
C8837 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00269f
C8838 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.79e-21
C8839 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 5.17e-21
C8840 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00305f
C8841 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 3.26e-21
C8842 sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__conb_1_15/HI 0.00406f
C8843 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_48/Y 0.0104f
C8844 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 5.33e-19
C8845 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0211f
C8846 sky130_fd_sc_hd__dfbbn_1_26/Q_N V_LOW -0.00253f
C8847 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 4.35e-20
C8848 sky130_fd_sc_hd__inv_16_20/A sky130_fd_sc_hd__inv_16_7/Y 1.28e-19
C8849 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# -0.00786f
C8850 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0.021f
C8851 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_647_21# 0.0025f
C8852 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# V_LOW 4.8e-20
C8853 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# -0.00141f
C8854 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# V_LOW -0.00121f
C8855 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.3e-19
C8856 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# V_LOW 1.79e-20
C8857 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00321f
C8858 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__inv_1_10/Y 3.92e-20
C8859 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_18/A 0.232f
C8860 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.96e-20
C8861 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__inv_16_40/Y 1.5e-19
C8862 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q -5.74e-21
C8863 sky130_fd_sc_hd__dfbbn_1_46/a_557_413# V_LOW 3.56e-20
C8864 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__conb_1_20/HI 0.0115f
C8865 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 3.72e-19
C8866 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0417f
C8867 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0285f
C8868 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.166f
C8869 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 2.43e-20
C8870 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_66/A 5.65e-20
C8871 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 5.59e-21
C8872 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.66e-21
C8873 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# 0.00359f
C8874 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_58/Y 2.2e-21
C8875 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0216f
C8876 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_1_13/Y 0.00313f
C8877 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# 0.00742f
C8878 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_16_41/Y 0.0317f
C8879 sky130_fd_sc_hd__dfbbn_1_16/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 5.22e-20
C8880 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.106f
C8881 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# -0.00889f
C8882 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 1.04e-19
C8883 sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__inv_1_14/Y 0.00391f
C8884 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 3.5e-19
C8885 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# V_LOW -0.00121f
C8886 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_51/Y 0.00349f
C8887 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# V_LOW -2.68e-19
C8888 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__nand3_1_2/Y 0.0264f
C8889 sky130_fd_sc_hd__fill_4_194/VPB V_LOW 0.797f
C8890 sky130_fd_sc_hd__conb_1_5/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0195f
C8891 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_43/HI 2.48e-20
C8892 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0317f
C8893 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.44e-19
C8894 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_24/HI 8.31e-20
C8895 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# sky130_fd_sc_hd__conb_1_44/HI 9.79e-19
C8896 sky130_fd_sc_hd__conb_1_28/LO RISING_COUNTER.COUNT_SUB_DFF10.Q 1.8e-20
C8897 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__conb_1_48/HI 3.24e-19
C8898 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00255f
C8899 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# V_LOW -0.0272f
C8900 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# -0.00385f
C8901 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# sky130_fd_sc_hd__inv_1_41/Y 6.02e-20
C8902 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1_24/LO 4.57e-20
C8903 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.016f
C8904 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0169f
C8905 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0396f
C8906 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 8.26e-20
C8907 FULL_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0141f
C8908 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0317f
C8909 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0834f
C8910 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 0.00113f
C8911 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.329f
C8912 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0433f
C8913 sky130_fd_sc_hd__inv_16_20/A sky130_fd_sc_hd__inv_1_67/A 0.00855f
C8914 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 1.97e-19
C8915 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 1.97e-19
C8916 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 5.81e-19
C8917 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.0167f
C8918 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.29e-19
C8919 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# V_LOW 0.00251f
C8920 sky130_fd_sc_hd__conb_1_7/LO RISING_COUNTER.COUNT_SUB_DFF8.Q 1.04e-19
C8921 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# -0.0496f
C8922 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# -2.65e-20
C8923 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 0.0035f
C8924 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 3.22e-20
C8925 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_29/Y 4.39e-22
C8926 sky130_fd_sc_hd__nand3_1_0/a_109_47# V_LOW -2.94e-19
C8927 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_581_47# -2.6e-20
C8928 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 9.79e-19
C8929 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__conb_1_47/HI 0.134f
C8930 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 6.76e-21
C8931 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 1.35e-20
C8932 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 1.49e-20
C8933 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_581_47# 2.86e-19
C8934 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 5.25e-20
C8935 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_29/A 0.0404f
C8936 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 6.36e-20
C8937 sky130_fd_sc_hd__conb_1_17/HI sky130_fd_sc_hd__conb_1_19/HI 3.29e-20
C8938 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_39/LO 1.7e-20
C8939 sky130_fd_sc_hd__dfbbn_1_44/Q_N RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0272f
C8940 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# V_LOW 0.00546f
C8941 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 8.07e-20
C8942 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 0.00106f
C8943 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 0.00122f
C8944 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 5.05e-19
C8945 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 4.66e-19
C8946 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_40/Y 0.92f
C8947 sky130_fd_sc_hd__conb_1_49/HI V_LOW 0.0657f
C8948 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_647_21# -6.43e-20
C8949 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_473_413# -3.06e-20
C8950 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# -0.00336f
C8951 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_381_47# -3.79e-20
C8952 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# sky130_fd_sc_hd__conb_1_20/HI 0.0176f
C8953 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.00691f
C8954 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# 9.5e-20
C8955 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0299f
C8956 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 0.026f
C8957 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.45e-19
C8958 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.45e-19
C8959 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0179f
C8960 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__conb_1_11/LO 5.27e-20
C8961 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.014f
C8962 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_64/A 5.63e-20
C8963 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_27/Y 0.0668f
C8964 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__nand3_1_1/Y 0.00209f
C8965 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00234f
C8966 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00462f
C8967 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__conb_1_24/HI 0.00481f
C8968 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 9.65e-21
C8969 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.51e-20
C8970 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1_7/HI 0.00153f
C8971 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/Q_N 4.32e-19
C8972 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_58/Y 6.25e-19
C8973 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0102f
C8974 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.0247f
C8975 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__nand2_1_2/A 2.37e-20
C8976 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# V_LOW 0.0139f
C8977 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__conb_1_50/HI 2.11e-20
C8978 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0405f
C8979 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_56/A 0.0114f
C8980 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_13/LO 7.28e-19
C8981 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__conb_1_9/HI 0.0143f
C8982 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_581_47# -2.6e-20
C8983 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0.00387f
C8984 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_30/HI 1.67e-20
C8985 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# -4.37e-20
C8986 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# -6.22e-19
C8987 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# -6.23e-21
C8988 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00108f
C8989 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00502f
C8990 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0121f
C8991 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_55/Y 0.0923f
C8992 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 1.89e-19
C8993 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__inv_1_39/Y 4.43e-21
C8994 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 9.19e-21
C8995 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0287f
C8996 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0431f
C8997 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_10/Y 0.00248f
C8998 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__conb_1_10/HI 0.0114f
C8999 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 2.89e-19
C9000 sky130_fd_sc_hd__fill_4_184/VPB V_LOW 0.797f
C9001 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# sky130_fd_sc_hd__conb_1_48/HI -0.00243f
C9002 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0557f
C9003 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# V_LOW -0.00251f
C9004 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.52e-20
C9005 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00661f
C9006 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 0.0049f
C9007 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 0.0388f
C9008 sky130_fd_sc_hd__conb_1_9/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.56e-20
C9009 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__nand2_8_8/A 0.0163f
C9010 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# 9.52e-19
C9011 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1_19/Y 4.48e-20
C9012 sky130_fd_sc_hd__inv_1_2/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 8.79e-20
C9013 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 1.58e-19
C9014 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_19/Y 0.00127f
C9015 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0634f
C9016 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 0.0125f
C9017 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_1_27/Y 5.25e-21
C9018 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# -0.00624f
C9019 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_557_413# -3.67e-20
C9020 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00201f
C9021 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# sky130_fd_sc_hd__inv_1_0/Y 0.00307f
C9022 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.38e-20
C9023 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_48/Y 8.88e-19
C9024 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__nor2_1_0/Y 1.04e-19
C9025 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_1_41/Y 0.146f
C9026 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 4.35e-21
C9027 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_7/A 0.151f
C9028 sky130_fd_sc_hd__conb_1_14/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 3.99e-19
C9029 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_26/Y 1.7e-19
C9030 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_18/A 2.53e-19
C9031 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 8.29e-20
C9032 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.00125f
C9033 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.108f
C9034 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00303f
C9035 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 2.38e-19
C9036 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 3.27e-19
C9037 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# V_LOW 2.03e-19
C9038 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_1_49/Y 0.248f
C9039 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0.0301f
C9040 sky130_fd_sc_hd__conb_1_46/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0314f
C9041 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# 4.17e-20
C9042 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00389f
C9043 sky130_fd_sc_hd__inv_1_34/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0637f
C9044 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 6.21e-20
C9045 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 2.93e-20
C9046 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_19/Q_N 0.03f
C9047 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# 3.12e-19
C9048 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_8_0/A 0.0038f
C9049 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0514f
C9050 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.21e-19
C9051 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__conb_1_51/HI 6.06e-19
C9052 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 0.00108f
C9053 sky130_fd_sc_hd__conb_1_13/HI FULL_COUNTER.COUNT_SUB_DFF17.Q 0.253f
C9054 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 1.39e-19
C9055 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 2.62e-19
C9056 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# sky130_fd_sc_hd__inv_1_26/Y 4.15e-20
C9057 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.0208f
C9058 sky130_fd_sc_hd__inv_1_35/Y V_LOW 0.131f
C9059 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__inv_1_2/Y 0.00318f
C9060 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# V_LOW 0.00407f
C9061 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_1_30/Y 6.44e-20
C9062 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 9.86e-20
C9063 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 4.77e-20
C9064 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0244f
C9065 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__inv_16_41/Y 6.49e-20
C9066 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# -5.54e-21
C9067 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -2.18e-19
C9068 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# -9.62e-19
C9069 sky130_fd_sc_hd__conb_1_4/HI FULL_COUNTER.COUNT_SUB_DFF6.Q 2.09e-20
C9070 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00493f
C9071 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__inv_1_24/Y 4.06e-20
C9072 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# sky130_fd_sc_hd__conb_1_50/HI -6.57e-19
C9073 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__conb_1_28/HI 3.76e-21
C9074 sky130_fd_sc_hd__inv_1_3/Y V_LOW 2.7f
C9075 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 3.33e-21
C9076 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# 3.49e-21
C9077 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__conb_1_3/HI 0.00947f
C9078 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 0.00145f
C9079 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__nand3_1_2/Y 0.00115f
C9080 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00103f
C9081 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__conb_1_2/HI 3.04e-21
C9082 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.13e-21
C9083 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_4_0/A 9.87e-20
C9084 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.006f
C9085 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.92e-20
C9086 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 5.5e-21
C9087 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_1_34/Y 1.31e-20
C9088 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.47e-19
C9089 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.153f
C9090 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_20/HI 9.87e-21
C9091 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# sky130_fd_sc_hd__conb_1_14/HI 0.0015f
C9092 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__conb_1_9/HI 0.00123f
C9093 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_1_63/Y 8.12e-22
C9094 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0361f
C9095 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__inv_1_35/Y 0.128f
C9096 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 1.43e-20
C9097 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 2.07e-20
C9098 sky130_fd_sc_hd__dfbbn_1_10/Q_N FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0312f
C9099 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 0.00192f
C9100 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__conb_1_39/HI 2e-19
C9101 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 3.26e-19
C9102 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# sky130_fd_sc_hd__inv_1_50/Y 1.05e-20
C9103 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__conb_1_32/HI 0.00472f
C9104 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.451f
C9105 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__conb_1_33/HI 1.18e-19
C9106 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_1_67/A 3.88e-19
C9107 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# Reset 0.00714f
C9108 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_23/HI 0.0204f
C9109 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# sky130_fd_sc_hd__inv_1_27/Y 7.69e-22
C9110 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 0.181f
C9111 sky130_fd_sc_hd__inv_16_9/A V_LOW 0.356f
C9112 FULL_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0304f
C9113 sky130_fd_sc_hd__nand2_8_1/a_27_47# V_LOW -0.0117f
C9114 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# -5.42e-19
C9115 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__inv_1_33/Y 2.33e-21
C9116 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.69e-20
C9117 sky130_fd_sc_hd__inv_16_16/Y sky130_fd_sc_hd__inv_16_15/A 0.0852f
C9118 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.00216f
C9119 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0147f
C9120 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__conb_1_2/HI 0.0261f
C9121 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_53/A 0.3f
C9122 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 4.88e-20
C9123 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# sky130_fd_sc_hd__inv_1_41/Y 0.00132f
C9124 sky130_fd_sc_hd__conb_1_11/HI V_LOW 0.0957f
C9125 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# sky130_fd_sc_hd__inv_1_59/Y 0.00162f
C9126 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.06e-21
C9127 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__conb_1_30/HI 4.84e-20
C9128 sky130_fd_sc_hd__nand2_1_2/A Reset 7.22e-19
C9129 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.69e-20
C9130 sky130_fd_sc_hd__inv_16_51/A sky130_fd_sc_hd__inv_16_50/A 0.00496f
C9131 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 8.3e-19
C9132 sky130_fd_sc_hd__conb_1_40/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.17e-19
C9133 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.28e-19
C9134 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# V_LOW 4.61e-20
C9135 sky130_fd_sc_hd__inv_16_22/A V_LOW 0.298f
C9136 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_39/HI 0.00127f
C9137 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# -0.00512f
C9138 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_557_413# -0.0012f
C9139 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__inv_1_1/Y 3.32e-20
C9140 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# -3.79e-20
C9141 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# -0.00336f
C9142 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 1.25e-19
C9143 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__inv_1_49/Y 0.00554f
C9144 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 6.53e-21
C9145 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_791_47# 0.00378f
C9146 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00148f
C9147 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00617f
C9148 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__inv_1_40/Y 0.101f
C9149 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00942f
C9150 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_65/Y 0.00395f
C9151 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# -1.67e-19
C9152 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# -0.00175f
C9153 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -6.22e-19
C9154 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_2_0/A 9.27e-20
C9155 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__inv_1_3/Y 1.07e-20
C9156 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.7e-21
C9157 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_2_0/A 0.00169f
C9158 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 0.00577f
C9159 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 1.97e-19
C9160 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.43e-20
C9161 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 9.92e-21
C9162 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.06e-20
C9163 sky130_fd_sc_hd__conb_1_3/LO FULL_COUNTER.COUNT_SUB_DFF7.Q 7.78e-21
C9164 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 0.0355f
C9165 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# sky130_fd_sc_hd__inv_1_2/Y 1.07e-21
C9166 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_66/A 0.00256f
C9167 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__inv_1_25/Y 6e-19
C9168 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.00211f
C9169 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# V_LOW -0.0978f
C9170 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# -9.32e-20
C9171 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# 2.84e-32
C9172 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -1.89e-19
C9173 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# -2.48e-19
C9174 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.82e-19
C9175 sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_9/Y 0.0767f
C9176 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.21e-19
C9177 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_1_60/Y 0.0262f
C9178 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__inv_1_50/Y 0.00262f
C9179 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/Q_N 0.00133f
C9180 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# -2.74e-21
C9181 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_66/A 0.0687f
C9182 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# V_LOW 2.26e-20
C9183 sky130_fd_sc_hd__conb_1_10/LO FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0171f
C9184 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 1.94e-21
C9185 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 6.97e-22
C9186 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 3.17e-19
C9187 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0387f
C9188 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0217f
C9189 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# 0.00123f
C9190 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_8_8/A 4.58e-19
C9191 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00277f
C9192 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_24/HI 2.26e-19
C9193 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_1_29/Y 0.0417f
C9194 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_56/A 0.0781f
C9195 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0.00139f
C9196 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 6.35e-19
C9197 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 5.67e-21
C9198 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1_36/Y 0.0434f
C9199 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00917f
C9200 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__conb_1_33/HI 3.25e-19
C9201 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_1_9/Y 8.62e-19
C9202 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_1/HI 0.0738f
C9203 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__inv_1_27/Y 0.0107f
C9204 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# Reset 2.16e-19
C9205 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# 0.00289f
C9206 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# CLOCK_GEN.SR_Op.Q 1.61e-19
C9207 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 0.0243f
C9208 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 4.29e-20
C9209 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 4.98e-21
C9210 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__inv_1_3/Y 2.73e-20
C9211 sky130_fd_sc_hd__conb_1_0/LO FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0413f
C9212 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_16/Y 0.0832f
C9213 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.22e-19
C9214 sky130_fd_sc_hd__nand2_8_2/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 6.21e-19
C9215 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__conb_1_33/LO 8.81e-20
C9216 RISING_COUNTER.COUNT_SUB_DFF4.Q V_LOW 1.46f
C9217 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_5/HI 0.0221f
C9218 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# sky130_fd_sc_hd__conb_1_29/HI 9.39e-20
C9219 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.81e-19
C9220 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -6.22e-19
C9221 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# -6.23e-21
C9222 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# -0.00175f
C9223 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# -0.00441f
C9224 FALLING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF9.Q 0.46f
C9225 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__inv_1_32/Y 0.0358f
C9226 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# 3.09e-19
C9227 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# V_LOW 0.0357f
C9228 sky130_fd_sc_hd__dfbbn_1_30/Q_N V_LOW -9.93e-19
C9229 sky130_fd_sc_hd__inv_1_63/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.36e-19
C9230 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__inv_1_41/Y 1.94e-20
C9231 RISING_COUNTER.COUNT_SUB_DFF1.Q Reset 0.0425f
C9232 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# -5.42e-19
C9233 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_8_0/A 0.0537f
C9234 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00169f
C9235 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 5.03e-20
C9236 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 5.09e-20
C9237 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.07e-19
C9238 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_66/Y 0.324f
C9239 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0.00382f
C9240 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 3.13e-19
C9241 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 0.00128f
C9242 RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00157f
C9243 FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00709f
C9244 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 3.01e-21
C9245 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__inv_1_38/Y 2.42e-19
C9246 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.00369f
C9247 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 7.3e-20
C9248 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.07e-19
C9249 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__conb_1_39/LO 0.0174f
C9250 sky130_fd_sc_hd__conb_1_47/LO sky130_fd_sc_hd__conb_1_49/LO 0.00241f
C9251 sky130_fd_sc_hd__inv_1_37/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 6.25e-21
C9252 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# V_LOW 0.0143f
C9253 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_36/Y 0.00209f
C9254 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__inv_1_25/Y 0.00142f
C9255 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_31/HI 0.00441f
C9256 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_557_413# -3.67e-20
C9257 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# -0.0313f
C9258 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00321f
C9259 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_1_32/Y 9.25e-19
C9260 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# V_LOW -9.15e-19
C9261 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# V_LOW -0.00389f
C9262 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF12.Q 4.88e-21
C9263 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# V_LOW -2.68e-19
C9264 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.254f
C9265 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/Q_N -4.33e-20
C9266 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# -1.76e-19
C9267 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__inv_1_59/Y 0.0155f
C9268 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# V_LOW 0.00509f
C9269 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 3.87e-19
C9270 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_25/LO 9.17e-19
C9271 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# -0.00794f
C9272 sky130_fd_sc_hd__dfbbn_1_23/Q_N FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.19e-19
C9273 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 2.86e-19
C9274 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# Reset 0.027f
C9275 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_47/Y 0.0104f
C9276 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_67/A 0.00176f
C9277 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_66/A 0.00961f
C9278 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__inv_16_40/Y 0.3f
C9279 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_1_44/A 0.283f
C9280 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_557_413# 0.00224f
C9281 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__conb_1_19/HI 1.68e-19
C9282 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# V_LOW 0.0185f
C9283 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 6.04e-20
C9284 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI 0.00337f
C9285 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 0.00231f
C9286 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.49e-19
C9287 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00291f
C9288 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__nor2_1_0/Y 0.0329f
C9289 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_36/LO 1.27e-20
C9290 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.4e-19
C9291 sky130_fd_sc_hd__conb_1_27/LO V_LOW 0.0988f
C9292 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 2.68e-19
C9293 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 2.68e-19
C9294 sky130_fd_sc_hd__conb_1_14/LO FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00205f
C9295 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__inv_1_60/Y 5.65e-19
C9296 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 8.4e-21
C9297 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 6.66e-19
C9298 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.003f
C9299 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 9.05e-19
C9300 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 1.86e-21
C9301 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 4.59e-19
C9302 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00169f
C9303 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_44/A 0.00176f
C9304 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_3/A 0.00733f
C9305 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.35e-20
C9306 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0685f
C9307 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__inv_1_43/Y 0.0466f
C9308 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# sky130_fd_sc_hd__inv_16_40/Y 0.00101f
C9309 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__conb_1_33/HI 0.00104f
C9310 sky130_fd_sc_hd__inv_1_19/Y V_LOW 0.188f
C9311 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__conb_1_37/HI 0.00984f
C9312 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.173f
C9313 sky130_fd_sc_hd__conb_1_38/LO V_LOW 0.0966f
C9314 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.0172f
C9315 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# V_LOW 0.00675f
C9316 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# CLOCK_GEN.SR_Op.Q 5.53e-20
C9317 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 9.5e-21
C9318 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 7.79e-20
C9319 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.94e-21
C9320 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_791_47# 0.00656f
C9321 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.53e-19
C9322 sky130_fd_sc_hd__inv_1_51/Y V_LOW 0.112f
C9323 sky130_fd_sc_hd__conb_1_16/LO V_LOW 0.0479f
C9324 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 1.16e-19
C9325 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 5.3e-19
C9326 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 2.14e-19
C9327 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__nand2_8_9/A 1.07e-20
C9328 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.81e-21
C9329 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 3.95e-19
C9330 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00201f
C9331 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# -0.00141f
C9332 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_1_38/Y 2.12e-21
C9333 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__nand2_1_2/A 0.00113f
C9334 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0427f
C9335 sky130_fd_sc_hd__dfbbn_1_42/Q_N FALLING_COUNTER.COUNT_SUB_DFF8.Q 8.03e-19
C9336 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# V_LOW 2.94e-20
C9337 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# sky130_fd_sc_hd__inv_1_28/Y 5.21e-19
C9338 V_SENSE sky130_fd_sc_hd__inv_16_6/A 0.78f
C9339 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_19/A 0.0998f
C9340 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_2_0/A 0.285f
C9341 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# 5.42e-20
C9342 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_31/HI 5.88e-20
C9343 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# V_LOW 0.014f
C9344 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_891_329# 0.00119f
C9345 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_65/Y 7.43e-20
C9346 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_8_0/Y 4.11e-19
C9347 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/Q_N -9.56e-20
C9348 sky130_fd_sc_hd__conb_1_9/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 4.01e-20
C9349 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_17/HI 7.02e-19
C9350 sky130_fd_sc_hd__inv_1_42/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0909f
C9351 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__inv_1_38/Y 4.71e-19
C9352 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.66e-19
C9353 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# 2.65e-19
C9354 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_30/Y 0.0416f
C9355 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# 1.24e-19
C9356 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__conb_1_29/LO 4.72e-20
C9357 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# -0.00497f
C9358 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# sky130_fd_sc_hd__inv_16_41/Y 3e-20
C9359 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0148f
C9360 sky130_fd_sc_hd__conb_1_45/LO FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00316f
C9361 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__inv_1_36/Y 1.64e-20
C9362 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 3.86e-20
C9363 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_35/Y 0.188f
C9364 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_66/A 0.0139f
C9365 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 6.16e-21
C9366 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 0.00217f
C9367 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00309f
C9368 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 1.71e-20
C9369 sky130_fd_sc_hd__dfbbn_1_49/a_581_47# sky130_fd_sc_hd__inv_1_59/Y 2.47e-19
C9370 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# V_LOW 0.0422f
C9371 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# V_LOW 1.57e-20
C9372 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_1_39/Y 0.00947f
C9373 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF15.Q 4.41e-21
C9374 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 8.34e-21
C9375 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_41/Y 0.0395f
C9376 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -7.6e-19
C9377 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# -5.54e-21
C9378 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__conb_1_16/HI 0.0346f
C9379 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_581_47# -2.6e-20
C9380 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# Reset 2.47e-19
C9381 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__inv_1_44/A 0.0011f
C9382 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/Q_N -4.24e-20
C9383 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_18/LO 9.45e-19
C9384 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_10/Y 0.247f
C9385 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# V_LOW 0.00451f
C9386 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 8.07e-21
C9387 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__inv_1_48/Y 1.16e-19
C9388 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__inv_1_7/Y 0.0061f
C9389 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.86e-19
C9390 FALLING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 9.87e-21
C9391 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# 3.97e-19
C9392 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# V_LOW 2.26e-20
C9393 sky130_fd_sc_hd__inv_1_36/Y V_LOW 0.0516f
C9394 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_17/Q_N 2.4e-19
C9395 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.00619f
C9396 sky130_fd_sc_hd__inv_1_34/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.36e-20
C9397 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/Q_N 0.011f
C9398 sky130_fd_sc_hd__conb_1_33/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0326f
C9399 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_381_47# -2.53e-20
C9400 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_20/HI 0.0772f
C9401 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 8.03e-21
C9402 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00241f
C9403 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_891_329# -2.2e-20
C9404 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -0.0166f
C9405 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# V_LOW 2.86e-20
C9406 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__conb_1_30/HI 0.00434f
C9407 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_26/HI 0.00181f
C9408 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.23e-19
C9409 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/Q_N 7.01e-20
C9410 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.15e-22
C9411 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 3.44e-21
C9412 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__conb_1_28/LO 1.67e-19
C9413 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0265f
C9414 sky130_fd_sc_hd__inv_16_19/Y V_LOW 0.185f
C9415 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# V_LOW 1.38e-19
C9416 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_17/LO 0.0471f
C9417 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0207f
C9418 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00442f
C9419 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 2.93e-20
C9420 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_1/Y 0.186f
C9421 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__inv_1_10/Y 0.00245f
C9422 sky130_fd_sc_hd__dfbbn_1_43/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0126f
C9423 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0162f
C9424 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__conb_1_42/LO 0.00206f
C9425 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_40/HI 2.04e-19
C9426 sky130_fd_sc_hd__inv_16_41/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.115f
C9427 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_34/LO 6.9e-19
C9428 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 0.887f
C9429 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# -1.46e-20
C9430 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# -0.00222f
C9431 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_47/Y 1.75e-19
C9432 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# V_LOW -0.116f
C9433 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_24/Y 0.00537f
C9434 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0247f
C9435 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 3.38e-20
C9436 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 0.0209f
C9437 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.07e-19
C9438 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# sky130_fd_sc_hd__conb_1_47/HI 6.14e-19
C9439 sky130_fd_sc_hd__inv_1_23/A V_LOW 0.329f
C9440 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0198f
C9441 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_29/LO 3.81e-20
C9442 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# -0.00141f
C9443 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# -0.00717f
C9444 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_557_413# -3.67e-20
C9445 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 5.87e-21
C9446 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__nand3_1_2/Y 2.5e-21
C9447 sky130_fd_sc_hd__conb_1_45/HI sky130_fd_sc_hd__inv_1_59/Y 0.0398f
C9448 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_2/Y 0.276f
C9449 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# V_LOW -1.01e-19
C9450 sky130_fd_sc_hd__dfbbn_1_32/Q_N V_LOW -5.13e-19
C9451 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00102f
C9452 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# -3.34e-20
C9453 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__conb_1_16/HI 0.00759f
C9454 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__inv_1_41/Y 0.0032f
C9455 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__conb_1_5/HI 1.58e-19
C9456 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__conb_1_18/LO 5.56e-19
C9457 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 8.78e-20
C9458 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 1.73e-19
C9459 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__conb_1_23/HI 0.016f
C9460 sky130_fd_sc_hd__conb_1_13/HI FULL_COUNTER.COUNT_SUB_DFF14.Q 7.43e-21
C9461 sky130_fd_sc_hd__nand2_8_8/A V_LOW 0.101f
C9462 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 8.78e-20
C9463 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# -1.44e-20
C9464 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 1.78e-21
C9465 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__conb_1_34/HI 0.00278f
C9466 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0091f
C9467 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 0.0901f
C9468 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__conb_1_20/HI 3.41e-19
C9469 sky130_fd_sc_hd__inv_1_40/Y V_LOW 0.221f
C9470 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 2.97e-19
C9471 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# 0.0012f
C9472 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_473_413# -0.0109f
C9473 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_647_21# -0.00631f
C9474 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__inv_1_37/Y 1.69e-20
C9475 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__inv_1_26/Y 2.86e-20
C9476 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00176f
C9477 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# -0.017f
C9478 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.326f
C9479 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# -0.00592f
C9480 sky130_fd_sc_hd__dfbbn_1_27/Q_N V_LOW -0.00128f
C9481 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__conb_1_13/HI 2.45e-19
C9482 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__conb_1_19/HI 5.57e-21
C9483 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__conb_1_30/HI 0.00139f
C9484 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 4.91e-20
C9485 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__inv_1_20/Y 6.92e-19
C9486 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.5e-19
C9487 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__inv_1_29/Y 1.75e-19
C9488 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 5.98e-19
C9489 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_34/LO 7.23e-20
C9490 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.00153f
C9491 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__conb_1_21/HI 1.22e-20
C9492 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.58e-20
C9493 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_1_31/Y 3.26e-20
C9494 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 3.75e-19
C9495 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00246f
C9496 sky130_fd_sc_hd__conb_1_51/LO FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0598f
C9497 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00242f
C9498 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 7.16e-20
C9499 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__inv_1_40/Y 0.00172f
C9500 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_24/HI 0.0104f
C9501 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_27/a_381_47# 4.51e-19
C9502 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 0.00122f
C9503 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 0.00122f
C9504 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__inv_1_38/Y 0.251f
C9505 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.37f
C9506 V_SENSE sky130_fd_sc_hd__inv_16_26/Y 1.43e-19
C9507 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.02e-19
C9508 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__conb_1_16/HI 3.35e-19
C9509 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/Q_N 2.11e-19
C9510 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 0.00542f
C9511 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# -9.32e-20
C9512 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 3.13e-19
C9513 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00382f
C9514 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 5.09e-20
C9515 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 0.00128f
C9516 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__inv_16_40/Y 8.21e-21
C9517 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# V_LOW -9.94e-19
C9518 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00341f
C9519 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 0.00114f
C9520 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/Q_N 0.00181f
C9521 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00313f
C9522 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__conb_1_25/HI 0.0115f
C9523 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# Reset 5.23e-20
C9524 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0024f
C9525 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_28/HI 1.35e-20
C9526 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_53/A 0.193f
C9527 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_66/Y 0.00127f
C9528 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__conb_1_17/HI 2.27e-20
C9529 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 8.43e-20
C9530 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 2.89e-21
C9531 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 9.93e-20
C9532 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 3.58e-20
C9533 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_25/Y 7.01e-20
C9534 sky130_fd_sc_hd__dfbbn_1_16/Q_N FULL_COUNTER.COUNT_SUB_DFF14.Q 3.96e-19
C9535 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# V_LOW 3.56e-20
C9536 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -0.00524f
C9537 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_891_329# -0.00159f
C9538 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__conb_1_4/HI 0.0116f
C9539 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.5e-19
C9540 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_50/HI 0.0916f
C9541 sky130_fd_sc_hd__conb_1_37/HI CLOCK_GEN.SR_Op.Q 0.0205f
C9542 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 4.41e-20
C9543 FALLING_COUNTER.COUNT_SUB_DFF3.Q V_LOW 1.15f
C9544 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/Q_N -4.78e-20
C9545 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0.00784f
C9546 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# sky130_fd_sc_hd__inv_1_41/Y 1.07e-21
C9547 sky130_fd_sc_hd__inv_16_28/Y V_LOW 0.334f
C9548 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.56e-19
C9549 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 2.03e-20
C9550 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 6.87e-20
C9551 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__conb_1_39/HI 3.76e-21
C9552 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -7.83e-20
C9553 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_473_413# -3.86e-20
C9554 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_45/Y 0.0272f
C9555 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_891_329# -0.00159f
C9556 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# -0.00882f
C9557 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# sky130_fd_sc_hd__conb_1_23/HI 1.26e-19
C9558 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_46/A 2.49e-19
C9559 sky130_fd_sc_hd__conb_1_28/LO RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00261f
C9560 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__inv_16_41/Y 0.0296f
C9561 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# V_LOW 0.0318f
C9562 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 6.87e-20
C9563 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.81e-19
C9564 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 0.00152f
C9565 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 5.37e-19
C9566 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 5.17e-20
C9567 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 2.96e-19
C9568 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00229f
C9569 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__inv_1_25/Y 0.0107f
C9570 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.34e-19
C9571 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__conb_1_20/HI 3.29e-20
C9572 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# sky130_fd_sc_hd__conb_1_38/HI 0.00138f
C9573 FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.161f
C9574 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_15/HI 5e-20
C9575 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 1.89e-20
C9576 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# V_LOW -0.069f
C9577 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# -1.27e-19
C9578 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 7.82e-19
C9579 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00127f
C9580 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.0345f
C9581 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_47/A 0.154f
C9582 sky130_fd_sc_hd__nand2_1_5/Y CLOCK_GEN.SR_Op.Q 5.46e-20
C9583 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__inv_1_3/Y 6.95e-21
C9584 sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# sky130_fd_sc_hd__conb_1_19/HI 4.08e-19
C9585 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__conb_1_30/HI -2.17e-19
C9586 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# sky130_fd_sc_hd__inv_1_34/Y 0.00135f
C9587 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF11.Q 1.79e-19
C9588 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 1.75e-19
C9589 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.00121f
C9590 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 5.12e-20
C9591 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.26f
C9592 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 9.26e-22
C9593 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# V_LOW 0.00577f
C9594 sky130_fd_sc_hd__conb_1_37/LO FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00436f
C9595 sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 2.14e-19
C9596 sky130_fd_sc_hd__dfbbn_1_5/Q_N FULL_COUNTER.COUNT_SUB_DFF12.Q 2.7e-20
C9597 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_39/LO 1.19e-20
C9598 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_10/HI 4.84e-20
C9599 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.129f
C9600 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# sky130_fd_sc_hd__conb_1_21/HI -4.57e-19
C9601 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.128f
C9602 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 0.00246f
C9603 V_HIGH RISING_COUNTER.COUNT_SUB_DFF4.Q 1.19f
C9604 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 3.75e-19
C9605 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_12/HI 0.0298f
C9606 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0.137f
C9607 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# sky130_fd_sc_hd__conb_1_24/HI -0.00262f
C9608 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__inv_1_38/Y 0.00727f
C9609 sky130_fd_sc_hd__nand2_8_7/a_27_47# CLOCK_GEN.SR_Op.Q 3.76e-19
C9610 sky130_fd_sc_hd__conb_1_45/HI sky130_fd_sc_hd__inv_1_58/Y 6.8e-19
C9611 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__conb_1_51/HI 4.28e-20
C9612 sky130_fd_sc_hd__inv_16_28/Y sky130_fd_sc_hd__inv_16_9/Y 0.0179f
C9613 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# Reset 1.05e-20
C9614 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.35e-20
C9615 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__conb_1_17/HI 0.00144f
C9616 sky130_fd_sc_hd__inv_8_0/Y V_LOW 0.158f
C9617 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# 2.02e-20
C9618 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/Q_N -4.24e-20
C9619 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# V_LOW 3.56e-20
C9620 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_10/HI 0.00244f
C9621 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.00114f
C9622 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 0.0116f
C9623 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 4.03e-19
C9624 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 0.0116f
C9625 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.00278f
C9626 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_29/HI -9.93e-19
C9627 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 1.51e-19
C9628 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.111f
C9629 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00291f
C9630 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.37e-20
C9631 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_51/Y 0.197f
C9632 sky130_fd_sc_hd__dfbbn_1_27/Q_N RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00109f
C9633 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00273f
C9634 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 4.72e-20
C9635 sky130_fd_sc_hd__dfbbn_1_21/Q_N FALLING_COUNTER.COUNT_SUB_DFF12.Q 8.59e-19
C9636 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 2.48e-19
C9637 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# sky130_fd_sc_hd__conb_1_25/HI 0.0176f
C9638 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.43e-21
C9639 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_44/HI 0.0354f
C9640 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 3.61e-20
C9641 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_43/HI 0.00542f
C9642 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_16_40/Y 1.6e-19
C9643 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_25/LO 1.03e-20
C9644 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# -2.3e-19
C9645 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_941_21# -3.07e-19
C9646 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 1.65e-19
C9647 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# Reset 0.0195f
C9648 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.083f
C9649 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.98e-20
C9650 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 4.56e-21
C9651 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# -0.00342f
C9652 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# -3.86e-20
C9653 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# -0.00385f
C9654 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.44e-20
C9655 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 0.102f
C9656 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 8.26e-21
C9657 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_581_47# 1.26e-19
C9658 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 7.67e-19
C9659 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 8.83e-19
C9660 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 5.03e-19
C9661 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# -0.00631f
C9662 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# -0.00988f
C9663 sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__inv_1_59/Y 0.00261f
C9664 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_24/A 4.36e-20
C9665 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 5e-19
C9666 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 8.64e-19
C9667 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# -2.57e-20
C9668 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__inv_1_31/Y 7.05e-20
C9669 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# -0.00385f
C9670 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -1.42e-32
C9671 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_32/HI 3.89e-21
C9672 sky130_fd_sc_hd__nand3_1_2/a_109_47# V_LOW -2.94e-19
C9673 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_381_47# 0.0112f
C9674 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 2.2e-20
C9675 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_381_47# 8.36e-19
C9676 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0273f
C9677 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# V_LOW 0.015f
C9678 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_56/A 0.00158f
C9679 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_791_47# 1.68e-19
C9680 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 5.22e-20
C9681 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 3.12e-20
C9682 sky130_fd_sc_hd__inv_16_6/A CLOCK_GEN.SR_Op.Q 2.83e-19
C9683 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_66/A 0.0285f
C9684 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 0.0123f
C9685 sky130_fd_sc_hd__conb_1_9/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 0.064f
C9686 sky130_fd_sc_hd__inv_16_23/A V_SENSE 0.00997f
C9687 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.164f
C9688 sky130_fd_sc_hd__inv_1_42/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 0.211f
C9689 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# -0.0179f
C9690 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.319f
C9691 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# V_LOW 0.0138f
C9692 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__conb_1_18/HI 0.00257f
C9693 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# V_LOW -2.68e-19
C9694 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/Q_N 0.0285f
C9695 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_581_47# -2.6e-20
C9696 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -0.0491f
C9697 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 0.127f
C9698 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.99e-19
C9699 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_14/HI 4.62e-19
C9700 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0106f
C9701 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# -0.00813f
C9702 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 6.42e-21
C9703 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00579f
C9704 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__conb_1_11/HI 1.98e-19
C9705 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_16_40/Y 0.00636f
C9706 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0652f
C9707 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0675f
C9708 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.0102f
C9709 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_29/Y 0.0747f
C9710 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# 2.48e-19
C9711 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# V_LOW -0.00389f
C9712 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# V_LOW -1.39e-35
C9713 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 3.58e-19
C9714 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_1_31/Y 3.98e-19
C9715 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 5.07e-19
C9716 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00214f
C9717 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.9e-22
C9718 sky130_fd_sc_hd__dfbbn_1_6/Q_N FULL_COUNTER.COUNT_SUB_DFF12.Q 6.44e-19
C9719 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 2.24e-19
C9720 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00176f
C9721 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__conb_1_12/HI 5.96e-19
C9722 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00609f
C9723 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__inv_1_37/Y 7.09e-19
C9724 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# Reset 7.29e-19
C9725 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# -4.66e-20
C9726 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_381_47# -3.79e-20
C9727 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# sky130_fd_sc_hd__conb_1_10/HI 0.00214f
C9728 sky130_fd_sc_hd__inv_1_47/Y V_LOW 0.612f
C9729 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.31e-19
C9730 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__conb_1_51/HI 0.0983f
C9731 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__conb_1_29/HI -3.88e-20
C9732 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0022f
C9733 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 5.2e-21
C9734 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00833f
C9735 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_1_2/A 0.0116f
C9736 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0031f
C9737 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__conb_1_26/HI 6.11e-20
C9738 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__conb_1_2/HI 2.24e-21
C9739 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 5.75e-20
C9740 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__dfbbn_1_26/Q_N 0.0284f
C9741 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__inv_1_50/Y 0.00648f
C9742 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__conb_1_50/HI 7.58e-19
C9743 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_16_42/Y 0.0228f
C9744 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# -0.00631f
C9745 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# sky130_fd_sc_hd__inv_1_33/Y 1.22e-21
C9746 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# -0.0109f
C9747 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__inv_16_41/Y 0.0127f
C9748 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# sky130_fd_sc_hd__conb_1_44/HI 5.29e-19
C9749 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00258f
C9750 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 8.95e-22
C9751 sky130_fd_sc_hd__inv_1_67/Y CLOCK_GEN.SR_Op.Q 0.102f
C9752 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# -1.65e-19
C9753 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# -7.17e-20
C9754 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.03f
C9755 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# Reset 0.00104f
C9756 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# -2.57e-20
C9757 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 3.54e-21
C9758 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# CLOCK_GEN.SR_Op.Q 0.00176f
C9759 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_16_2/Y 0.282f
C9760 sky130_fd_sc_hd__conb_1_29/HI V_LOW 0.0369f
C9761 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.1e-19
C9762 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00131f
C9763 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.0176f
C9764 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__conb_1_12/HI 0.00414f
C9765 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 1.61e-20
C9766 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__inv_16_41/Y 2.26e-20
C9767 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00131f
C9768 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00513f
C9769 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 0.00616f
C9770 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 1.9e-19
C9771 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__conb_1_3/HI 2.03e-19
C9772 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_43/LO 9.82e-19
C9773 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/Q_N -6.48e-19
C9774 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q -2.92e-20
C9775 sky130_fd_sc_hd__inv_16_41/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0388f
C9776 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.0231f
C9777 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_1_36/Y 8.34e-20
C9778 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# 8.91e-20
C9779 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 1.38e-20
C9780 RISING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 6f
C9781 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# -1.89e-19
C9782 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# -3.72e-19
C9783 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__conb_1_16/HI 8.67e-20
C9784 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 0.0209f
C9785 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__inv_1_12/Y 1.64e-20
C9786 V_SENSE sky130_fd_sc_hd__inv_16_32/Y 0.00123f
C9787 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.11e-20
C9788 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 0.00213f
C9789 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# V_LOW 2.26e-20
C9790 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# V_LOW 5.62e-20
C9791 V_SENSE sky130_fd_sc_hd__inv_1_60/Y 6.36e-19
C9792 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# sky130_fd_sc_hd__conb_1_18/HI 0.00163f
C9793 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0365f
C9794 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# V_LOW 3.56e-20
C9795 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.0445f
C9796 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_40/Y 2.97e-21
C9797 V_SENSE sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# 9.74e-20
C9798 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_24/Y 3.14e-21
C9799 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_26/HI 1.69e-19
C9800 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_21/LO 1.45e-19
C9801 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 0.165f
C9802 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_647_21# -0.00122f
C9803 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_473_413# -0.00312f
C9804 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 5.87e-20
C9805 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# -0.00107f
C9806 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00584f
C9807 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# V_LOW 1.38e-19
C9808 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 3.61e-19
C9809 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# sky130_fd_sc_hd__conb_1_11/HI -2.65e-20
C9810 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0154f
C9811 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.075f
C9812 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0423f
C9813 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 3.49e-19
C9814 sky130_fd_sc_hd__dfbbn_1_28/Q_N V_LOW 1.99e-19
C9815 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_67/A 1.45e-19
C9816 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_38/Y 2.11e-21
C9817 V_SENSE sky130_fd_sc_hd__fill_4_188/VPB 0.0211f
C9818 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_7/HI 4.42e-19
C9819 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.21e-19
C9820 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/Q_N 7.19e-19
C9821 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.2e-20
C9822 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_66/Y 1.41e-19
C9823 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0025f
C9824 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.0024f
C9825 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_1_44/A 0.0101f
C9826 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF7.Q 6.07e-19
C9827 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__inv_1_37/Y 1.58e-19
C9828 sky130_fd_sc_hd__inv_1_60/Y sky130_fd_sc_hd__inv_16_41/Y 1.34e-20
C9829 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_56/A 0.00141f
C9830 sky130_fd_sc_hd__dfbbn_1_47/Q_N Reset 0.00106f
C9831 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# V_LOW 3.56e-20
C9832 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# 8.67e-19
C9833 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 0.00136f
C9834 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 4.17e-20
C9835 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0.00384f
C9836 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# -6.23e-21
C9837 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# -3.03e-19
C9838 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.39e-20
C9839 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__conb_1_25/HI 0.00306f
C9840 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.00227f
C9841 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16_55/Y 0.045f
C9842 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_1_45/Y 2.77e-20
C9843 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.17e-19
C9844 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__conb_1_35/HI 2.66e-20
C9845 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_15/HI 6.84e-21
C9846 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.36e-19
C9847 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00523f
C9848 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__conb_1_12/HI 6.01e-21
C9849 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# sky130_fd_sc_hd__conb_1_50/HI 1.87e-20
C9850 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 7.05e-20
C9851 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# V_LOW 0.0127f
C9852 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.69e-19
C9853 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 0.00761f
C9854 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 7.18e-19
C9855 FALLING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 2.07f
C9856 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# V_LOW 3.53e-20
C9857 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00159f
C9858 sky130_fd_sc_hd__conb_1_33/LO RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00436f
C9859 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.7e-20
C9860 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 0.0105f
C9861 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 4.74e-20
C9862 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 7.23e-19
C9863 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 3.95e-19
C9864 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__conb_1_2/HI 1.45e-19
C9865 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_49/Y 1.33e-19
C9866 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00337f
C9867 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.00352f
C9868 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/Q_N 5.44e-19
C9869 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.41e-19
C9870 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00361f
C9871 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00606f
C9872 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# -0.00262f
C9873 sky130_fd_sc_hd__conb_1_10/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 0.074f
C9874 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__nor2_1_0/Y 4.78e-19
C9875 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 4.3e-21
C9876 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_2/Y 6.29e-19
C9877 sky130_fd_sc_hd__inv_1_53/Y Reset 2.42e-19
C9878 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# V_LOW 0.0165f
C9879 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__conb_1_33/HI 0.00879f
C9880 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_891_329# 0.00136f
C9881 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_12/HI 4.97e-19
C9882 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0221f
C9883 sky130_fd_sc_hd__dfbbn_1_1/a_581_47# sky130_fd_sc_hd__inv_16_40/Y 0.00217f
C9884 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0376f
C9885 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.129f
C9886 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# -1.66e-19
C9887 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 0.142f
C9888 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# -0.00263f
C9889 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__conb_1_31/HI -0.00233f
C9890 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_69/Y 0.0194f
C9891 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__conb_1_16/HI 1.69e-19
C9892 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_38/LO 0.00155f
C9893 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 0.00127f
C9894 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# -4.66e-20
C9895 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 1.67e-21
C9896 sky130_fd_sc_hd__dfbbn_1_31/Q_N V_LOW -9.22e-19
C9897 FALLING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 0.4f
C9898 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00686f
C9899 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0404f
C9900 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# V_LOW 0.0129f
C9901 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# sky130_fd_sc_hd__inv_16_40/Y 9.47e-19
C9902 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.0162f
C9903 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 9.31e-20
C9904 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_28/HI -0.00907f
C9905 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__conb_1_5/HI 4.95e-19
C9906 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__inv_1_32/Y 0.00992f
C9907 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_39/Y 1.31e-19
C9908 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00478f
C9909 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00558f
C9910 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__inv_1_25/Y 6.99e-19
C9911 sky130_fd_sc_hd__nand2_8_4/a_27_47# V_LOW -0.0051f
C9912 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# 0.00355f
C9913 sky130_fd_sc_hd__dfbbn_1_16/Q_N FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0156f
C9914 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__conb_1_0/HI 7.57e-21
C9915 FULL_COUNTER.COUNT_SUB_DFF8.Q V_LOW 1.55f
C9916 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__conb_1_32/HI 0.00176f
C9917 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_46/A 1.46e-19
C9918 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00334f
C9919 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.00401f
C9920 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 3.88e-19
C9921 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 9.08e-19
C9922 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 3.22e-19
C9923 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__conb_1_20/HI 9.39e-21
C9924 V_SENSE sky130_fd_sc_hd__fill_4_182/VPB 0.0211f
C9925 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0197f
C9926 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# sky130_fd_sc_hd__inv_1_44/A 0.0035f
C9927 sky130_fd_sc_hd__inv_1_63/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q 6.58e-21
C9928 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# 1.31e-20
C9929 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_3/HI 2.76e-21
C9930 RISING_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 3.59e-20
C9931 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 3.78e-19
C9932 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 2.12e-21
C9933 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_30/HI 0.00561f
C9934 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 1.07e-19
C9935 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.0161f
C9936 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_64/A 0.00275f
C9937 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_45/Y 1.3e-20
C9938 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# 1.52e-19
C9939 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.16e-19
C9940 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00153f
C9941 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__conb_1_0/HI 2.38e-19
C9942 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_59/Y 0.00282f
C9943 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# V_LOW 2.26e-20
C9944 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 0.018f
C9945 sky130_fd_sc_hd__conb_1_2/LO V_LOW 0.129f
C9946 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00109f
C9947 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# V_LOW 1.79e-20
C9948 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 2.92e-20
C9949 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0192f
C9950 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_24/Y 6.82e-20
C9951 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 4.74e-21
C9952 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_55/A 0.00355f
C9953 sky130_fd_sc_hd__dfbbn_1_5/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00185f
C9954 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_66/A 7.95e-20
C9955 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 6.48e-20
C9956 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.0303f
C9957 sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 2.6e-20
C9958 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.011f
C9959 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0447f
C9960 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 8.6e-19
C9961 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/Q_N 4.46e-21
C9962 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.0176f
C9963 sky130_fd_sc_hd__dfbbn_1_7/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00672f
C9964 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_6/HI 0.00261f
C9965 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# V_LOW 0.00599f
C9966 V_HIGH FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.567f
C9967 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 7.17e-21
C9968 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# -0.00108f
C9969 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_941_21# 0.0153f
C9970 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.18e-19
C9971 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0706f
C9972 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# -9.32e-20
C9973 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# sky130_fd_sc_hd__conb_1_31/HI -0.00261f
C9974 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__conb_1_16/HI 3e-19
C9975 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__inv_1_0/Y 1.51e-19
C9976 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00407f
C9977 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_15/HI 2.15e-19
C9978 sky130_fd_sc_hd__inv_16_20/A V_LOW 0.31f
C9979 sky130_fd_sc_hd__dfbbn_1_8/Q_N FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0198f
C9980 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q -4.43e-21
C9981 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_1_42/Y 0.0154f
C9982 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# -6.23e-21
C9983 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -8.96e-20
C9984 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_381_47# -4.37e-20
C9985 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__conb_1_28/HI -9.71e-19
C9986 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 2.78e-21
C9987 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 1.67e-21
C9988 sky130_fd_sc_hd__inv_16_49/A sky130_fd_sc_hd__inv_16_48/A 1.7f
C9989 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_1_60/Y 7.48e-20
C9990 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0216f
C9991 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_17/Q_N 0.0288f
C9992 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 7.32e-20
C9993 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 6e-21
C9994 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__conb_1_19/LO 1.22e-19
C9995 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__conb_1_2/HI 0.00114f
C9996 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 5.7e-19
C9997 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.85e-19
C9998 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00102f
C9999 sky130_fd_sc_hd__inv_1_48/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00807f
C10000 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.00485f
C10001 sky130_fd_sc_hd__dfbbn_1_46/Q_N FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.43e-19
C10002 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__inv_1_36/Y 0.00198f
C10003 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 3.29e-20
C10004 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# V_LOW 0.02f
C10005 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__conb_1_19/HI 1.29e-21
C10006 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# Reset 0.0179f
C10007 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0143f
C10008 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_33/Y 2.83e-20
C10009 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# -3.79e-20
C10010 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# -0.00336f
C10011 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00115f
C10012 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00501f
C10013 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 7.47e-19
C10014 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# -0.00393f
C10015 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_557_413# -0.0012f
C10016 sky130_fd_sc_hd__dfbbn_1_33/Q_N RISING_COUNTER.COUNT_SUB_DFF6.Q 5.13e-20
C10017 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_60/Y 0.273f
C10018 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# sky130_fd_sc_hd__conb_1_30/HI 5.75e-19
C10019 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 5.36e-22
C10020 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 1.45e-19
C10021 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_14/Y 0.0622f
C10022 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_16_40/Y 0.00318f
C10023 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# sky130_fd_sc_hd__conb_1_0/HI 4.32e-20
C10024 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0119f
C10025 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# sky130_fd_sc_hd__inv_1_31/Y 2.33e-20
C10026 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__conb_1_45/HI 0.00252f
C10027 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand2_8_9/A 6.97e-21
C10028 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.0286f
C10029 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0558f
C10030 sky130_fd_sc_hd__inv_1_66/A FULL_COUNTER.COUNT_SUB_DFF1.Q 1.31e-20
C10031 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00127f
C10032 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.51e-20
C10033 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__nor2_1_0/Y 3.05e-21
C10034 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 8.9e-21
C10035 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 5.16e-20
C10036 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_49/A 0.0207f
C10037 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/Q_N 1.97e-21
C10038 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.39e-19
C10039 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_32/Y 1.47e-19
C10040 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand3_1_1/Y 0.0733f
C10041 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_29/HI 1.18e-20
C10042 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# sky130_fd_sc_hd__inv_1_10/Y 2.91e-19
C10043 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__conb_1_50/HI 3.15e-19
C10044 FULL_COUNTER.COUNT_SUB_DFF2.Q transmission_gate_9/GN 0.108f
C10045 sky130_fd_sc_hd__nand2_8_2/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00164f
C10046 sky130_fd_sc_hd__dfbbn_1_6/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0304f
C10047 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/a_647_21# 4.15e-21
C10048 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# V_LOW -1.39e-35
C10049 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 1.22e-20
C10050 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 7.89e-19
C10051 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 3.92e-19
C10052 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 1.99e-19
C10053 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.74e-20
C10054 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_581_47# -2.6e-20
C10055 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# 2.5e-21
C10056 sky130_fd_sc_hd__inv_1_34/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 3.98e-20
C10057 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__inv_1_28/Y 0.00648f
C10058 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__inv_16_40/Y 1.86e-19
C10059 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__inv_2_0/A 0.0313f
C10060 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_16_40/Y 0.0327f
C10061 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__conb_1_7/HI 1.2e-21
C10062 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/Q_N -4.78e-20
C10063 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_1_21/Y 0.00183f
C10064 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.1e-19
C10065 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/Q_N 9.65e-21
C10066 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_13/HI 0.00886f
C10067 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# -1.69e-19
C10068 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 0.0455f
C10069 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.35e-20
C10070 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_16_40/Y 0.609f
C10071 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_49/A 5.49e-19
C10072 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__conb_1_17/HI 0.0223f
C10073 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__conb_1_28/HI -2.17e-19
C10074 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 6.89e-19
C10075 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00917f
C10076 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 1.59e-20
C10077 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__inv_1_60/Y 1.5e-19
C10078 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.301f
C10079 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 7.27e-20
C10080 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 8.14e-21
C10081 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand2_8_1/a_27_47# 8.88e-20
C10082 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 2.2e-20
C10083 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# sky130_fd_sc_hd__conb_1_2/HI 3.29e-20
C10084 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# V_LOW 1.38e-19
C10085 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_29/Y 1.02e-19
C10086 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_58/Y 0.105f
C10087 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 4.85e-19
C10088 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# 0.00178f
C10089 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# Reset 0.00409f
C10090 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0111f
C10091 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# CLOCK_GEN.SR_Op.Q 0.11f
C10092 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# V_LOW 0.00669f
C10093 sky130_fd_sc_hd__inv_16_41/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.119f
C10094 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 0.326f
C10095 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 6.53e-20
C10096 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__inv_1_1/Y 3.75e-21
C10097 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.09e-21
C10098 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0354f
C10099 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__conb_1_6/HI 0.0586f
C10100 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# 2.39e-19
C10101 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 8.46e-21
C10102 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.02e-19
C10103 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__inv_1_60/Y 5.46e-19
C10104 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# -0.0306f
C10105 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_557_413# -3.67e-20
C10106 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 2.2e-19
C10107 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0616f
C10108 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.25e-20
C10109 sky130_fd_sc_hd__inv_1_63/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0181f
C10110 sky130_fd_sc_hd__dfbbn_1_17/a_557_413# V_LOW 3.56e-20
C10111 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_1_39/Y -0.0038f
C10112 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__inv_16_40/Y 6.16e-19
C10113 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0761f
C10114 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.0263f
C10115 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 0.0168f
C10116 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.104f
C10117 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# 3.26e-19
C10118 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_47/Y 5.84e-19
C10119 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_61/Y 0.0381f
C10120 Reset sky130_fd_sc_hd__inv_1_49/Y 2.46e-20
C10121 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__conb_1_4/HI 4.08e-19
C10122 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 9.46e-20
C10123 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_16_40/Y 0.148f
C10124 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 7.8e-21
C10125 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__inv_1_38/Y 0.00953f
C10126 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_29/HI 8.03e-19
C10127 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__inv_1_32/Y 3.01e-19
C10128 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.81e-21
C10129 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__conb_1_26/HI -9.62e-19
C10130 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# -0.00381f
C10131 sky130_fd_sc_hd__dfbbn_1_45/Q_N V_LOW -0.00461f
C10132 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 5.58e-21
C10133 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__inv_1_27/Y 0.00324f
C10134 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00114f
C10135 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 2.08e-19
C10136 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 0.367f
C10137 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.11e-21
C10138 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_15/LO 0.0543f
C10139 V_SENSE sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 1.84e-20
C10140 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_44/A 0.00502f
C10141 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_4_0/A 3.49e-20
C10142 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0855f
C10143 sky130_fd_sc_hd__inv_1_60/Y sky130_fd_sc_hd__inv_1_63/Y 0.00446f
C10144 sky130_fd_sc_hd__inv_16_7/A V_LOW 0.0993f
C10145 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_581_47# -7.91e-19
C10146 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__inv_1_41/Y 0.132f
C10147 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_1_3/a_113_47# 5.84e-19
C10148 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_1_29/Y 3.56e-20
C10149 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_49/Y 2.17e-19
C10150 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__conb_1_15/HI 7.45e-20
C10151 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.282f
C10152 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# -4.66e-20
C10153 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# -3.79e-20
C10154 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/Q_N 9.65e-21
C10155 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.292f
C10156 sky130_fd_sc_hd__conb_1_33/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.23e-20
C10157 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# sky130_fd_sc_hd__inv_1_55/Y 0.00136f
C10158 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF17.Q 2.51e-20
C10159 sky130_fd_sc_hd__conb_1_22/LO FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0278f
C10160 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__conb_1_15/HI 0.0187f
C10161 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_2/Y 1.49e-20
C10162 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0504f
C10163 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 6.83e-20
C10164 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00152f
C10165 sky130_fd_sc_hd__conb_1_4/HI V_LOW 0.165f
C10166 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 7.67e-19
C10167 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# -0.00511f
C10168 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# V_LOW 0.0385f
C10169 sky130_fd_sc_hd__dfbbn_1_35/Q_N Reset 0.0166f
C10170 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# V_LOW -9.15e-19
C10171 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 4.84e-20
C10172 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_22/a_381_47# 1.16e-20
C10173 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# CLOCK_GEN.SR_Op.Q 0.0269f
C10174 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# -0.028f
C10175 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_557_413# -3.67e-20
C10176 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.76e-21
C10177 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# V_LOW -9.15e-19
C10178 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.11e-19
C10179 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# V_LOW 0.0194f
C10180 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_1_40/Y 6.07e-20
C10181 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__inv_1_11/Y 0.00134f
C10182 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__conb_1_7/HI 0.0192f
C10183 sky130_fd_sc_hd__nand2_8_2/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.85e-21
C10184 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 0.00189f
C10185 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0167f
C10186 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__conb_1_37/HI 1.59e-20
C10187 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# V_LOW -0.107f
C10188 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# V_LOW -0.00121f
C10189 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_38/HI 0.00328f
C10190 V_SENSE sky130_fd_sc_hd__inv_16_23/Y 0.00164f
C10191 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__inv_1_8/Y 7.11e-19
C10192 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 1.97e-21
C10193 sky130_fd_sc_hd__conb_1_26/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.56e-20
C10194 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__conb_1_4/HI 5.86e-21
C10195 RISING_COUNTER.COUNT_SUB_DFF3.Q V_LOW 1.35f
C10196 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_29/LO 1.7e-20
C10197 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__conb_1_24/HI 0.0482f
C10198 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_53/A 0.306f
C10199 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00126f
C10200 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 3.22e-20
C10201 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__inv_1_62/Y 4.44e-20
C10202 V_SENSE sky130_fd_sc_hd__inv_16_3/A 0.0544f
C10203 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# -1.44e-20
C10204 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# V_LOW 0.0134f
C10205 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 6.21e-19
C10206 sky130_fd_sc_hd__inv_1_56/Y CLOCK_GEN.SR_Op.Q 8.95e-19
C10207 sky130_fd_sc_hd__inv_16_42/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 0.11f
C10208 FULL_COUNTER.COUNT_SUB_DFF15.Q V_LOW 2.33f
C10209 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__conb_1_44/HI 0.0336f
C10210 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_2_0/A 0.016f
C10211 V_SENSE RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0384f
C10212 FALLING_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 1.2e-20
C10213 FULL_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 2.05e-19
C10214 RISING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.023f
C10215 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# -3.79e-20
C10216 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# -4.66e-20
C10217 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__inv_1_41/Y 7.08e-21
C10218 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00433f
C10219 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__inv_1_44/A 0.00288f
C10220 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 4.56e-20
C10221 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# V_LOW -0.00371f
C10222 sky130_fd_sc_hd__inv_1_50/Y V_LOW 0.399f
C10223 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__conb_1_8/LO 0.0127f
C10224 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.25e-19
C10225 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_19/Y 7.92e-20
C10226 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_39/HI 4.26e-21
C10227 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.25e-19
C10228 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00223f
C10229 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.78e-19
C10230 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.6e-21
C10231 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0407f
C10232 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 6.51e-20
C10233 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00414f
C10234 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 1.49e-20
C10235 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# sky130_fd_sc_hd__conb_1_15/HI -1.64e-20
C10236 sky130_fd_sc_hd__nand2_8_5/a_27_47# V_LOW -0.0117f
C10237 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.82e-20
C10238 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/Q_N 1.4e-20
C10239 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 1.81e-19
C10240 sky130_fd_sc_hd__nand3_1_0/Y Reset 0.0025f
C10241 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# sky130_fd_sc_hd__conb_1_8/HI 0.00138f
C10242 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_1_67/A 1.63e-20
C10243 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 3.14e-19
C10244 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 2.31e-19
C10245 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# -0.0105f
C10246 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# -0.00423f
C10247 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 0.00899f
C10248 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_581_47# -7.91e-19
C10249 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_16_41/Y 0.0311f
C10250 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# V_LOW 2.94e-20
C10251 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_473_413# 0.00316f
C10252 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_17/HI 2.03e-19
C10253 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# -5.42e-19
C10254 sky130_fd_sc_hd__dfbbn_1_51/Q_N V_LOW 1.99e-19
C10255 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# V_LOW -0.00266f
C10256 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_16_4/Y 1.67e-20
C10257 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.48e-19
C10258 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_14/LO 8.63e-20
C10259 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# V_LOW 0.011f
C10260 sky130_fd_sc_hd__dfbbn_1_13/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0232f
C10261 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_193_47# -0.0253f
C10262 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 3.47e-19
C10263 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 9.38e-21
C10264 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 2.42e-20
C10265 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__nand3_1_1/Y 0.00552f
C10266 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__conb_1_7/HI -6.37e-19
C10267 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00633f
C10268 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 8.12e-22
C10269 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__conb_1_31/HI 0.00103f
C10270 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# V_LOW 2.26e-20
C10271 RISING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 7.29e-19
C10272 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_557_413# 7.19e-19
C10273 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 0.00115f
C10274 sky130_fd_sc_hd__conb_1_51/HI Reset 0.0827f
C10275 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0193f
C10276 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__nand2_8_4/Y 3.26e-19
C10277 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# V_LOW -9.94e-19
C10278 sky130_fd_sc_hd__inv_16_6/A FALLING_COUNTER.COUNT_SUB_DFF4.Q 7.11e-20
C10279 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0868f
C10280 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 1.71e-20
C10281 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_24/HI 0.0281f
C10282 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.022f
C10283 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.59e-21
C10284 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# 7.12e-19
C10285 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_58/Y 3.35e-21
C10286 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0274f
C10287 sky130_fd_sc_hd__nor2_1_0/Y V_LOW 0.304f
C10288 sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__inv_1_40/Y 0.00767f
C10289 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# -0.00431f
C10290 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# -0.00458f
C10291 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0317f
C10292 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.72e-19
C10293 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# V_LOW -0.00266f
C10294 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__inv_1_69/Y 5.2e-20
C10295 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# V_LOW 0.0117f
C10296 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_16_42/Y 0.0267f
C10297 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__conb_1_40/HI 0.00126f
C10298 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__conb_1_43/HI 1.49e-20
C10299 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0356f
C10300 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.237f
C10301 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_24/HI 1.42e-19
C10302 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_4_0/A 0.122f
C10303 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# sky130_fd_sc_hd__conb_1_44/HI 6.75e-19
C10304 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0032f
C10305 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# V_LOW -0.00809f
C10306 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__conb_1_48/HI 0.0328f
C10307 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 5.85e-20
C10308 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00525f
C10309 sky130_fd_sc_hd__inv_1_2/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0222f
C10310 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.72e-19
C10311 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 2.45e-19
C10312 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.6e-20
C10313 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_1_44/A 2.09e-19
C10314 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 2.82e-20
C10315 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.0181f
C10316 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0201f
C10317 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00814f
C10318 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 0.0272f
C10319 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.35e-20
C10320 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0459f
C10321 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.48e-19
C10322 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00209f
C10323 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_31/HI 1.83e-19
C10324 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 0.32f
C10325 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.334f
C10326 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# V_LOW -2.84e-19
C10327 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0164f
C10328 sky130_fd_sc_hd__inv_1_64/A V_LOW -0.00461f
C10329 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# -1.27e-19
C10330 sky130_fd_sc_hd__inv_1_65/A FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00347f
C10331 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.83e-20
C10332 sky130_fd_sc_hd__nand3_1_0/a_193_47# V_LOW -5.03e-19
C10333 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# 0.00534f
C10334 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_16_19/Y 0.00189f
C10335 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__conb_1_12/HI 0.00202f
C10336 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 0.347f
C10337 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__conb_1_40/HI -0.00465f
C10338 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# sky130_fd_sc_hd__conb_1_17/HI 9.65e-21
C10339 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__nand2_8_0/a_27_47# 6.28e-19
C10340 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00138f
C10341 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.12e-19
C10342 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 5.29e-21
C10343 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# V_LOW 0.0133f
C10344 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 0.0035f
C10345 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 0.0029f
C10346 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 0.00106f
C10347 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_941_21# -0.00409f
C10348 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_473_413# -3.86e-20
C10349 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 6.6e-19
C10350 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__nand3_1_1/Y 0.0678f
C10351 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 0.0351f
C10352 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.00666f
C10353 sky130_fd_sc_hd__conb_1_22/HI FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.01e-19
C10354 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.42e-20
C10355 sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# sky130_fd_sc_hd__conb_1_20/HI -2.65e-20
C10356 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00216f
C10357 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.99e-19
C10358 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 1.99e-19
C10359 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.19e-19
C10360 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.19e-19
C10361 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0317f
C10362 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_47/A 5.27e-19
C10363 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_47/A 4.4e-20
C10364 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.036f
C10365 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00888f
C10366 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# sky130_fd_sc_hd__conb_1_24/HI 5.29e-19
C10367 sky130_fd_sc_hd__conb_1_5/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0103f
C10368 sky130_fd_sc_hd__conb_1_1/LO V_LOW 0.0499f
C10369 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__conb_1_20/HI 0.0116f
C10370 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_36/LO 0.0116f
C10371 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00402f
C10372 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.6e-19
C10373 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 3.01e-20
C10374 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__nand2_1_2/A 1.63e-20
C10375 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.00556f
C10376 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.0604f
C10377 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.23e-20
C10378 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# V_LOW 0.0153f
C10379 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0748f
C10380 sky130_fd_sc_hd__conb_1_24/HI V_LOW 0.169f
C10381 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_47/Q_N 0.00266f
C10382 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_13/LO 5.9e-20
C10383 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__conb_1_9/HI 0.0107f
C10384 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0.00103f
C10385 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__conb_1_20/HI 9.65e-19
C10386 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0361f
C10387 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# -2.53e-20
C10388 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00272f
C10389 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 6.78e-20
C10390 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 4.96e-20
C10391 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__inv_1_39/Y 1.87e-20
C10392 V_SENSE RISING_COUNTER.COUNT_SUB_DFF1.Q 6.43e-20
C10393 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_6/Y 2.93e-19
C10394 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_13/LO 6.57e-20
C10395 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0297f
C10396 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0402f
C10397 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00196f
C10398 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_14/HI 0.0352f
C10399 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_10/HI 7.45e-20
C10400 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_3/Y 3e-19
C10401 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand2_8_8/A 0.262f
C10402 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# sky130_fd_sc_hd__conb_1_48/HI 7e-19
C10403 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0194f
C10404 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 7.23e-21
C10405 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__conb_1_39/HI 8.76e-19
C10406 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 6.12e-20
C10407 sky130_fd_sc_hd__dfbbn_1_29/Q_N RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0296f
C10408 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 0.0446f
C10409 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 0.0219f
C10410 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 0.002f
C10411 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 0.0353f
C10412 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_16_4/Y 0.00234f
C10413 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__inv_1_9/Y 5.95e-22
C10414 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF16.Q 6.94e-19
C10415 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00764f
C10416 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_891_329# 0.00134f
C10417 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__inv_1_27/Y 1.59e-19
C10418 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_891_329# -2.2e-20
C10419 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# -9.65e-20
C10420 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.25e-19
C10421 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__conb_1_31/HI 3.29e-20
C10422 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# sky130_fd_sc_hd__inv_1_0/Y 4.53e-19
C10423 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 3.44e-20
C10424 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 8.87e-20
C10425 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__inv_1_12/Y 2.27e-20
C10426 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_41/Y 0.223f
C10427 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_44/A 0.0562f
C10428 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__inv_1_62/Y 0.0145f
C10429 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_25/LO 2.56e-19
C10430 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_581_47# -2.6e-20
C10431 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_1_31/Y 6.68e-19
C10432 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_1_41/Y 0.0972f
C10433 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_66/A 0.346f
C10434 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.35e-19
C10435 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_46/Q_N 0.00148f
C10436 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 4.38e-21
C10437 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 3.28e-21
C10438 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 2.06e-20
C10439 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 9.09e-22
C10440 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 1.18e-21
C10441 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.048f
C10442 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.91e-19
C10443 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# V_LOW 1.38e-19
C10444 sky130_fd_sc_hd__conb_1_31/HI V_LOW 0.126f
C10445 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# V_LOW 1.79e-20
C10446 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# -0.0139f
C10447 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__inv_1_49/Y 0.0256f
C10448 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 0.0162f
C10449 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# 5.74e-20
C10450 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# -9.41e-19
C10451 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00386f
C10452 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_11/HI 0.389f
C10453 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# 0.00164f
C10454 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0.00136f
C10455 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.00384f
C10456 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 4.17e-20
C10457 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 8.67e-19
C10458 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 2.1e-19
C10459 sky130_fd_sc_hd__nand3_1_2/Y V_LOW 1.29f
C10460 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0397f
C10461 sky130_fd_sc_hd__conb_1_3/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 0.135f
C10462 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.56e-19
C10463 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_0/a_27_47# 8e-19
C10464 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__conb_1_51/HI 3.28e-19
C10465 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# 0.00987f
C10466 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 1.99e-20
C10467 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 0.00784f
C10468 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__inv_1_26/Y 2.55e-19
C10469 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.0143f
C10470 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.034f
C10471 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00207f
C10472 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__inv_1_2/Y 1.72e-20
C10473 sky130_fd_sc_hd__inv_1_54/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.143f
C10474 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# V_LOW 0.00433f
C10475 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 1.14e-20
C10476 sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# sky130_fd_sc_hd__inv_16_41/Y 3.64e-19
C10477 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# -1.67e-19
C10478 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -9.88e-20
C10479 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# -0.00175f
C10480 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16_48/A 0.00154f
C10481 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_31/HI 1e-19
C10482 sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# sky130_fd_sc_hd__conb_1_9/HI -8.7e-21
C10483 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 0.00733f
C10484 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__conb_1_3/HI 0.00492f
C10485 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# -1.44e-20
C10486 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 5.44e-19
C10487 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_16_8/A 6.59e-21
C10488 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__nand3_1_2/Y 5.84e-19
C10489 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0034f
C10490 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_21/Y 0.00359f
C10491 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_49/Y 0.0091f
C10492 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.87e-21
C10493 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__conb_1_8/HI 9.56e-19
C10494 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 4.84e-21
C10495 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00635f
C10496 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.03e-19
C10497 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 7.1e-20
C10498 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 4.75e-21
C10499 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__inv_1_34/Y 0.0108f
C10500 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0631f
C10501 sky130_fd_sc_hd__dfbbn_1_11/Q_N FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0237f
C10502 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# sky130_fd_sc_hd__conb_1_14/HI 1.57e-19
C10503 sky130_fd_sc_hd__conb_1_48/HI RISING_COUNTER.COUNT_SUB_DFF9.Q 0.037f
C10504 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 0.00282f
C10505 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_9/HI 0.00141f
C10506 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.01e-20
C10507 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.53e-19
C10508 sky130_fd_sc_hd__dfbbn_1_36/Q_N V_LOW -0.00993f
C10509 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__inv_1_63/Y 9.58e-21
C10510 sky130_fd_sc_hd__dfbbn_1_31/a_581_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00217f
C10511 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_473_413# 5.62e-19
C10512 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__conb_1_39/HI 1.3e-19
C10513 sky130_fd_sc_hd__conb_1_9/HI V_LOW 0.176f
C10514 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0432f
C10515 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__nand2_8_8/A 5.15e-19
C10516 sky130_fd_sc_hd__dfbbn_1_13/Q_N FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0233f
C10517 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# Reset 0.00341f
C10518 sky130_fd_sc_hd__conb_1_0/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 1.05e-20
C10519 sky130_fd_sc_hd__conb_1_24/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0267f
C10520 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_23/HI 0.0228f
C10521 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_2_0/A 9.87e-21
C10522 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__inv_1_27/Y 3.87e-19
C10523 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0.113f
C10524 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# -0.00282f
C10525 sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0141f
C10526 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 0.00144f
C10527 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.00201f
C10528 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.74e-20
C10529 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 7.48e-20
C10530 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00452f
C10531 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__conb_1_2/HI 0.00942f
C10532 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.79e-20
C10533 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__inv_1_41/Y 0.0388f
C10534 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__inv_1_59/Y 0.00307f
C10535 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 2.67e-20
C10536 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__conb_1_29/HI 6.79e-20
C10537 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_2_0/A 0.0883f
C10538 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_52/A 0.186f
C10539 sky130_fd_sc_hd__inv_1_40/Y sky130_fd_sc_hd__inv_1_38/Y 3.01e-21
C10540 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 7.48e-20
C10541 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 8.65e-19
C10542 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.022f
C10543 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00265f
C10544 sky130_fd_sc_hd__inv_1_2/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00115f
C10545 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 6.66e-20
C10546 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__inv_1_1/Y 7.53e-21
C10547 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# -0.00524f
C10548 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_891_329# -0.00159f
C10549 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.75e-20
C10550 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# sky130_fd_sc_hd__inv_1_49/Y 6.07e-19
C10551 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 3.96e-19
C10552 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0268f
C10553 RISING_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.925f
C10554 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__inv_1_40/Y 7.91e-19
C10555 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__inv_1_35/Y 0.00108f
C10556 sky130_fd_sc_hd__inv_16_40/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0288f
C10557 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 3.78e-19
C10558 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0173f
C10559 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# -0.00441f
C10560 sky130_fd_sc_hd__fill_8_958/VPB V_LOW 0.797f
C10561 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_47/A 0.0271f
C10562 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_2_0/A 2.21e-19
C10563 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0155f
C10564 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__inv_1_3/Y 0.00843f
C10565 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_40/a_27_47# 1.72e-19
C10566 sky130_fd_sc_hd__conb_1_46/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0306f
C10567 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 1.21e-19
C10568 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00342f
C10569 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# 2.53e-19
C10570 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 0.0123f
C10571 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 4.99e-19
C10572 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 2.23e-20
C10573 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.73e-21
C10574 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 0.00182f
C10575 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.81e-20
C10576 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_64/Y 3.41e-20
C10577 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# V_LOW 1.79e-20
C10578 sky130_fd_sc_hd__conb_1_7/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 1.52e-20
C10579 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 6.29e-19
C10580 sky130_fd_sc_hd__dfbbn_1_5/Q_N FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00882f
C10581 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_52/A 0.105f
C10582 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# V_LOW 0.0177f
C10583 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_3/HI 2.1e-20
C10584 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# -2.74e-21
C10585 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -2.18e-19
C10586 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# -1.6e-19
C10587 sky130_fd_sc_hd__conb_1_20/HI V_LOW 0.171f
C10588 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_19/A 0.321f
C10589 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00201f
C10590 sky130_fd_sc_hd__inv_16_2/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0852f
C10591 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# sky130_fd_sc_hd__conb_1_3/HI -0.00262f
C10592 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_1_60/Y 0.00312f
C10593 V_HIGH RISING_COUNTER.COUNT_SUB_DFF3.Q 1.49f
C10594 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_381_47# -3.04e-19
C10595 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# -6.23e-21
C10596 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__conb_1_41/LO 6.65e-19
C10597 sky130_fd_sc_hd__conb_1_23/LO V_LOW 0.0848f
C10598 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# V_LOW 4.8e-20
C10599 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 0.0156f
C10600 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.28e-20
C10601 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 1.28e-19
C10602 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 1.37e-20
C10603 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_28/Y 0.0623f
C10604 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00238f
C10605 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.0261f
C10606 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0497f
C10607 sky130_fd_sc_hd__inv_1_57/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 2.72e-20
C10608 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.23e-20
C10609 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.00152f
C10610 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 5.48e-21
C10611 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_1_29/Y 0.0566f
C10612 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# 5.88e-20
C10613 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 1.74e-20
C10614 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.4e-20
C10615 sky130_fd_sc_hd__conb_1_45/LO V_LOW 0.0518f
C10616 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_47/Y 3.1e-20
C10617 RISING_COUNTER.COUNT_SUB_DFF15.Q V_LOW 2.21f
C10618 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_1_9/Y 0.00102f
C10619 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# sky130_fd_sc_hd__inv_1_27/Y 8.17e-19
C10620 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# Reset 1.15e-20
C10621 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__conb_1_23/HI 0.00388f
C10622 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 0.0468f
C10623 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# CLOCK_GEN.SR_Op.Q 2.96e-19
C10624 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0276f
C10625 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_647_21# 0.0157f
C10626 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 0.00132f
C10627 sky130_fd_sc_hd__conb_1_34/LO V_LOW 0.0674f
C10628 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 4.22e-19
C10629 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__conb_1_2/HI -2.07e-19
C10630 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_17/HI 9.22e-20
C10631 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# -0.00441f
C10632 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# -0.0244f
C10633 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_557_413# -3.67e-20
C10634 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_15/A 0.102f
C10635 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_47/Y 0.00529f
C10636 sky130_fd_sc_hd__nand2_1_2/A CLOCK_GEN.SR_Op.Q 1.26e-19
C10637 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_37/HI 4.88e-19
C10638 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__inv_1_32/Y 0.00844f
C10639 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/Q_N 8.53e-21
C10640 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__conb_1_15/HI 1.36e-20
C10641 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# V_LOW 0.0204f
C10642 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_17/HI 0.127f
C10643 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# -0.00385f
C10644 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_52/A 0.00262f
C10645 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand3_1_2/a_193_47# 6.69e-20
C10646 sky130_fd_sc_hd__dfbbn_1_33/Q_N RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00187f
C10647 sky130_fd_sc_hd__conb_1_22/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 2.31e-19
C10648 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__inv_16_40/Y 9.92e-20
C10649 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_1/Y 8.2e-20
C10650 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00119f
C10651 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 0.00378f
C10652 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00347f
C10653 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# -0.00141f
C10654 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 0.00138f
C10655 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 9.2e-20
C10656 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00545f
C10657 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 1.98e-19
C10658 sky130_fd_sc_hd__conb_1_47/LO FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00292f
C10659 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_2_0/A 1.7e-21
C10660 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0472f
C10661 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_47/Y 0.13f
C10662 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 9.55e-19
C10663 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_34/LO 0.0523f
C10664 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__inv_1_38/Y 2.34e-21
C10665 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 3.95e-19
C10666 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# 2.32e-19
C10667 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_39/LO 6.66e-19
C10668 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 0.374f
C10669 sky130_fd_sc_hd__conb_1_44/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 2.47e-20
C10670 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__inv_1_36/Y 7.7e-21
C10671 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# V_LOW 0.0125f
C10672 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__conb_1_31/HI 1.18e-20
C10673 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 8.59e-20
C10674 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_891_329# -2.2e-20
C10675 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# -0.0139f
C10676 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__inv_1_32/Y 4.45e-19
C10677 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_66/A 0.0541f
C10678 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 3.81e-19
C10679 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# V_LOW -9.15e-19
C10680 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# V_LOW -0.00121f
C10681 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 9.42e-21
C10682 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_35/Y 1.06e-19
C10683 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# V_LOW 0.00532f
C10684 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_30/Y 1.45e-20
C10685 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.101f
C10686 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# -9.32e-20
C10687 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/Q_N -9.56e-20
C10688 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__inv_1_59/Y 0.0167f
C10689 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# V_LOW 1.38e-19
C10690 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.17f
C10691 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# -0.00431f
C10692 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# -0.0105f
C10693 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__conb_1_28/HI 0.00329f
C10694 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF17.Q 0.004f
C10695 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# Reset 0.0267f
C10696 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_1_44/A 0.111f
C10697 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_891_329# 0.00295f
C10698 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 3.54e-21
C10699 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00309f
C10700 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# V_LOW 0.00585f
C10701 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 1.29e-19
C10702 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 9e-19
C10703 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 4.14e-21
C10704 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00493f
C10705 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__nor2_1_0/Y 0.00184f
C10706 sky130_fd_sc_hd__conb_1_3/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.92e-20
C10707 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00483f
C10708 sky130_fd_sc_hd__inv_16_32/Y sky130_fd_sc_hd__inv_16_8/A 0.00744f
C10709 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.59e-19
C10710 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__conb_1_7/LO 0.00256f
C10711 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 1.74e-19
C10712 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 1.74e-19
C10713 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 0.0256f
C10714 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 1.99e-20
C10715 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 1.99e-20
C10716 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__conb_1_15/HI 5.64e-21
C10717 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.0116f
C10718 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00278f
C10719 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 0.0116f
C10720 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 4.03e-19
C10721 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.00114f
C10722 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# sky130_fd_sc_hd__inv_1_29/Y 1.26e-20
C10723 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 8.26e-21
C10724 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_49/Y 2.7e-20
C10725 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00269f
C10726 sky130_fd_sc_hd__inv_16_27/Y sky130_fd_sc_hd__inv_16_29/Y 0.189f
C10727 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 4.95e-20
C10728 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_1_43/Y 0.0149f
C10729 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.119f
C10730 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__conb_1_37/HI 0.00294f
C10731 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_55/Y 0.242f
C10732 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_2/Y 0.0565f
C10733 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 0.0012f
C10734 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__conb_1_37/HI 2.26e-19
C10735 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0953f
C10736 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0351f
C10737 sky130_fd_sc_hd__conb_1_29/LO RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00578f
C10738 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 1.83e-20
C10739 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# V_LOW 1.38e-19
C10740 sky130_fd_sc_hd__inv_1_65/Y V_LOW 0.0248f
C10741 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.3e-20
C10742 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 9.72e-20
C10743 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.66e-19
C10744 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.0337f
C10745 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.0134f
C10746 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_581_47# 1.83e-19
C10747 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 1.73e-20
C10748 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 3.46e-20
C10749 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.23e-20
C10750 sky130_fd_sc_hd__inv_1_60/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.11e-21
C10751 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 0.00451f
C10752 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.00417f
C10753 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 3.14e-20
C10754 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.93e-20
C10755 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_49/Y 0.16f
C10756 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# -1.44e-20
C10757 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 7.53e-20
C10758 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# sky130_fd_sc_hd__inv_1_32/Y 2.05e-21
C10759 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0358f
C10760 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# sky130_fd_sc_hd__inv_1_28/Y 9.76e-19
C10761 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# V_LOW 4.73e-19
C10762 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/Q_N -6.48e-19
C10763 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_39/Y 1.05e-19
C10764 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__nand2_1_5/Y 0.0044f
C10765 sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 4.04e-20
C10766 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_31/HI 5.38e-21
C10767 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# V_LOW 0.0112f
C10768 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0288f
C10769 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# 8e-21
C10770 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__dfbbn_1_31/a_193_47# 3.67e-21
C10771 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 6.51e-20
C10772 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# 0.00417f
C10773 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__inv_1_1/Y 5.09e-21
C10774 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0077f
C10775 sky130_fd_sc_hd__conb_1_50/HI V_LOW 0.117f
C10776 sky130_fd_sc_hd__dfbbn_1_29/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.18e-19
C10777 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__inv_1_14/Y 0.0878f
C10778 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_17/HI 2.9e-19
C10779 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00176f
C10780 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_30/Y 0.0304f
C10781 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_8/A 1.22e-19
C10782 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_557_413# -3.67e-20
C10783 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# -0.0306f
C10784 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00215f
C10785 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__conb_1_31/HI 2.71e-21
C10786 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# -0.00592f
C10787 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 2.26e-21
C10788 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_1_35/Y 0.00602f
C10789 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 0.0287f
C10790 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.00336f
C10791 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/Q_N -4.78e-20
C10792 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0415f
C10793 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# V_LOW -0.309f
C10794 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.93e-20
C10795 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_1_39/Y 1.54e-19
C10796 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.00133f
C10797 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__conb_1_16/HI 0.00184f
C10798 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -6.22e-19
C10799 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# -6.23e-21
C10800 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# -0.00538f
C10801 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__inv_1_44/A 0.0199f
C10802 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# V_LOW 7.67e-22
C10803 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# V_LOW 4.8e-20
C10804 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.23e-19
C10805 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.56e-19
C10806 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_557_413# -3.67e-20
C10807 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_891_329# -2.46e-19
C10808 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# -5.33e-20
C10809 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 1.34e-19
C10810 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 1.34e-19
C10811 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 0.0185f
C10812 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.66e-19
C10813 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# sky130_fd_sc_hd__inv_1_43/Y 2.5e-21
C10814 sky130_fd_sc_hd__conb_1_42/LO V_LOW 0.0962f
C10815 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__conb_1_41/HI 0.0882f
C10816 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# sky130_fd_sc_hd__conb_1_41/HI 0.00212f
C10817 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0944f
C10818 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0391f
C10819 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# -4.66e-20
C10820 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# -3.79e-20
C10821 sky130_fd_sc_hd__inv_1_66/Y V_LOW 0.226f
C10822 sky130_fd_sc_hd__conb_1_33/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0183f
C10823 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__conb_1_30/HI 1.22e-20
C10824 V_SENSE sky130_fd_sc_hd__conb_1_44/HI 4.83e-19
C10825 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_16_4/Y 1.86e-20
C10826 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_44/Y 0.209f
C10827 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0548f
C10828 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# V_LOW 3.56e-20
C10829 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 5.7e-19
C10830 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0158f
C10831 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0224f
C10832 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 7.01e-20
C10833 sky130_fd_sc_hd__conb_1_35/HI V_LOW 0.0154f
C10834 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00386f
C10835 transmission_gate_9/GN FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.146f
C10836 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_40/HI 9.64e-20
C10837 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_31/HI 1.82e-20
C10838 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# -0.00216f
C10839 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# -0.00367f
C10840 V_SENSE sky130_fd_sc_hd__inv_16_24/Y 0.0279f
C10841 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__conb_1_17/HI 0.00154f
C10842 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# V_LOW -0.0245f
C10843 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_16_41/Y 2.87e-20
C10844 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0156f
C10845 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# sky130_fd_sc_hd__conb_1_47/HI 0.00211f
C10846 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_1_38/Y 1.39e-19
C10847 FULL_COUNTER.COUNT_SUB_DFF3.Q V_LOW 0.874f
C10848 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_891_329# -2.2e-20
C10849 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# -0.00953f
C10850 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 1.04e-19
C10851 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_1_35/Y 3.77e-20
C10852 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 7.22e-19
C10853 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__nand3_1_2/Y 2.55e-20
C10854 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__conb_1_40/HI 0.00365f
C10855 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_12/HI 0.0335f
C10856 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 6.53e-19
C10857 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__inv_1_39/Y 2.09e-19
C10858 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF15.Q 1.25e-19
C10859 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__conb_1_16/HI 0.00355f
C10860 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_1_41/Y 9.78e-20
C10861 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 1.13e-21
C10862 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# sky130_fd_sc_hd__conb_1_8/HI 9.74e-19
C10863 sky130_fd_sc_hd__dfbbn_1_24/Q_N V_LOW -0.00509f
C10864 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__conb_1_23/HI 0.00561f
C10865 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_34/Q_N 5.1e-20
C10866 FALLING_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 4.11f
C10867 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 2.77e-19
C10868 sky130_fd_sc_hd__inv_16_40/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0242f
C10869 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_17/HI -7.06e-21
C10870 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# sky130_fd_sc_hd__conb_1_34/HI 3.78e-19
C10871 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_38/HI 0.0108f
C10872 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0258f
C10873 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0325f
C10874 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__conb_1_27/HI 0.0301f
C10875 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__conb_1_20/HI 0.00306f
C10876 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF13.Q 5.04e-21
C10877 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_67/A 3.7e-20
C10878 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_381_47# 1.5e-21
C10879 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_1_45/Y 0.0132f
C10880 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_473_413# -0.0103f
C10881 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_941_21# -4.94e-19
C10882 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_1_48/Y 0.0167f
C10883 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0176f
C10884 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0249f
C10885 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# -1.27e-19
C10886 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0198f
C10887 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_16_4/Y 0.114f
C10888 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF12.Q 1.7e-19
C10889 sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# sky130_fd_sc_hd__conb_1_30/HI 3.38e-19
C10890 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.00885f
C10891 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.74e-19
C10892 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_2/HI 3.41e-20
C10893 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_34/LO 1.97e-35
C10894 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.00858f
C10895 sky130_fd_sc_hd__inv_16_2/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 2.23f
C10896 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_47/Y 0.071f
C10897 sky130_fd_sc_hd__conb_1_38/LO Reset 5.1e-21
C10898 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00413f
C10899 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0195f
C10900 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__conb_1_17/HI 1.75e-20
C10901 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__conb_1_38/HI 0.0025f
C10902 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.69e-20
C10903 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.48e-19
C10904 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 0.00275f
C10905 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_27/a_557_413# 9.05e-20
C10906 sky130_fd_sc_hd__inv_1_51/Y Reset 0.00177f
C10907 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 0.0048f
C10908 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__inv_1_38/Y 0.0264f
C10909 sky130_fd_sc_hd__inv_1_52/Y V_LOW 0.00431f
C10910 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__conb_1_16/HI 1.96e-20
C10911 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__nand2_8_8/A 1.22e-21
C10912 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0.0074f
C10913 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0.00138f
C10914 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 9.2e-20
C10915 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 1.98e-19
C10916 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.00545f
C10917 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 0.00378f
C10918 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# V_LOW -0.0125f
C10919 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.48e-19
C10920 V_SENSE sky130_fd_sc_hd__inv_16_47/Y 0.371f
C10921 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00137f
C10922 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 2.48e-19
C10923 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# -0.00592f
C10924 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_56/A 0.0531f
C10925 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# Reset 3.38e-20
C10926 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.43e-19
C10927 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.87e-19
C10928 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__inv_1_35/Y 6.2e-20
C10929 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# sky130_fd_sc_hd__conb_1_12/HI 0.00189f
C10930 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# V_LOW 2.26e-20
C10931 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# -0.00336f
C10932 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__conb_1_4/HI 0.00492f
C10933 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.21e-19
C10934 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 1.33e-19
C10935 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_17/HI 0.156f
C10936 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.00107f
C10937 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00612f
C10938 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__conb_1_16/HI 0.0233f
C10939 sky130_fd_sc_hd__fill_4_320/VPB V_LOW 0.797f
C10940 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__inv_1_58/Y 0.0135f
C10941 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.23e-19
C10942 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# -2.52e-19
C10943 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -4.72e-20
C10944 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# sky130_fd_sc_hd__conb_1_23/HI 0.00206f
C10945 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# -0.00336f
C10946 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# -3.79e-20
C10947 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# V_LOW 0.00352f
C10948 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# sky130_fd_sc_hd__conb_1_17/HI -2.22e-20
C10949 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__nand2_8_1/a_27_47# 8.06e-20
C10950 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0037f
C10951 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 5.61e-20
C10952 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 2.35e-19
C10953 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 2.16e-19
C10954 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 3.19e-21
C10955 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 3.41e-19
C10956 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 5.16e-19
C10957 sky130_fd_sc_hd__dfbbn_1_17/a_557_413# sky130_fd_sc_hd__inv_1_25/Y 8.17e-19
C10958 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__conb_1_27/HI -0.0127f
C10959 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 7.06e-21
C10960 RISING_COUNTER.COUNT_SUB_DFF0.Q transmission_gate_9/GN 0.0734f
C10961 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# V_LOW 0.026f
C10962 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0573f
C10963 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_5/A 7.26e-19
C10964 sky130_fd_sc_hd__inv_1_9/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 3.74e-21
C10965 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# -6.8e-19
C10966 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# -0.00631f
C10967 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# -0.00591f
C10968 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0317f
C10969 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_581_47# -2.6e-20
C10970 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00637f
C10971 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__inv_1_7/Y 3.69e-20
C10972 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0353f
C10973 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_16_4/Y 0.645f
C10974 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 1.44e-19
C10975 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0336f
C10976 FALLING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.743f
C10977 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_16_4/Y 1.25e-19
C10978 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 1.11e-20
C10979 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# V_LOW 1.38e-19
C10980 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 2.88e-20
C10981 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_66/A 1.83e-20
C10982 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__conb_1_34/LO 5.78e-20
C10983 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_39/LO 8.82e-19
C10984 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__inv_16_41/Y 8.09e-19
C10985 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__conb_1_10/HI 2.67e-20
C10986 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.078f
C10987 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_1_10/Y 1.63e-20
C10988 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0114f
C10989 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__conb_1_51/HI 2.54e-19
C10990 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__conb_1_12/HI 0.0173f
C10991 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 0.146f
C10992 sky130_fd_sc_hd__dfbbn_1_50/a_581_47# sky130_fd_sc_hd__inv_1_38/Y 6.07e-19
C10993 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.00472f
C10994 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__conb_1_5/HI 6.79e-20
C10995 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__nand2_8_4/Y 2.68e-20
C10996 sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__inv_1_66/Y 8.44e-21
C10997 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# Reset 4.52e-20
C10998 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_193_47# -0.135f
C10999 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 0.0594f
C11000 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# V_LOW 2.26e-20
C11001 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__conb_1_10/HI 0.0431f
C11002 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/Q_N -9.56e-20
C11003 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0502f
C11004 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 7.34e-19
C11005 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 9.14e-19
C11006 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 1e-19
C11007 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.001f
C11008 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__conb_1_29/HI -1.56e-20
C11009 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00127f
C11010 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 8.32e-19
C11011 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 9.75e-21
C11012 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.48e-21
C11013 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__conb_1_26/HI 7.33e-20
C11014 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__conb_1_31/HI 1.77e-19
C11015 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_46/A 0.00722f
C11016 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# sky130_fd_sc_hd__conb_1_25/HI -2.65e-20
C11017 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 0.0061f
C11018 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_27/Y 0.0196f
C11019 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.82e-20
C11020 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 0.0277f
C11021 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__conb_1_43/HI 0.00307f
C11022 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# -0.00263f
C11023 sky130_fd_sc_hd__inv_16_49/A sky130_fd_sc_hd__inv_16_50/A 3.34f
C11024 sky130_fd_sc_hd__inv_16_51/Y sky130_fd_sc_hd__inv_16_48/A 0.135f
C11025 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 2.2e-20
C11026 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0354f
C11027 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_47/Y 8.87e-20
C11028 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# Reset 0.0117f
C11029 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__nand2_8_4/Y 4.99e-19
C11030 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 2.84e-32
C11031 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_25/LO 5.37e-20
C11032 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.89e-19
C11033 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# -8.01e-19
C11034 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# -0.0014f
C11035 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__inv_1_9/Y 0.00234f
C11036 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# sky130_fd_sc_hd__conb_1_4/HI -0.00257f
C11037 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 0.0295f
C11038 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.54e-19
C11039 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_24/Y 1.16e-19
C11040 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00107f
C11041 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# 0.00156f
C11042 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.0123f
C11043 RISING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.28e-20
C11044 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# -0.0103f
C11045 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# -4.98e-19
C11046 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.2e-19
C11047 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 3.79e-20
C11048 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.54e-19
C11049 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# -1.76e-19
C11050 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_791_47# -2.22e-34
C11051 sky130_fd_sc_hd__nand3_1_2/a_193_47# V_LOW -5.03e-19
C11052 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 1.67e-21
C11053 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/Q_N 3.79e-20
C11054 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0025f
C11055 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0177f
C11056 sky130_fd_sc_hd__dfbbn_1_29/Q_N RISING_COUNTER.COUNT_SUB_DFF5.Q 1.41e-19
C11057 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_791_47# 9.9e-20
C11058 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 2.09e-19
C11059 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__inv_1_12/Y 5.19e-21
C11060 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# -1.69e-19
C11061 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0728f
C11062 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 0.406f
C11063 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# V_LOW 1.38e-19
C11064 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__conb_1_46/HI 0.00878f
C11065 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__conb_1_18/HI 6.77e-19
C11066 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# V_LOW 0.00994f
C11067 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_3/Y 0.0266f
C11068 sky130_fd_sc_hd__nand2_8_8/A Reset 0.0049f
C11069 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_44/A 8.37e-21
C11070 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# -6.78e-19
C11071 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_36/LO 7.17e-21
C11072 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 0.135f
C11073 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__conb_1_14/HI 1.75e-19
C11074 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# sky130_fd_sc_hd__inv_1_7/Y 2.32e-20
C11075 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00812f
C11076 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_557_413# -0.0012f
C11077 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# -0.00335f
C11078 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.36e-20
C11079 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.81e-19
C11080 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 2.58e-20
C11081 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 4.48e-21
C11082 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0378f
C11083 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.00265f
C11084 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# V_LOW -9.15e-19
C11085 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_51/Y 1.25f
C11086 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 1.31e-19
C11087 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 7.75e-22
C11088 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_44/HI 3.26e-20
C11089 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0194f
C11090 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.1e-21
C11091 sky130_fd_sc_hd__inv_16_29/A sky130_fd_sc_hd__inv_16_8/Y 0.0905f
C11092 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 3.73e-20
C11093 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.29e-19
C11094 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00859f
C11095 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__conb_1_14/HI 1.83e-20
C11096 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_1_30/Y 1.17e-19
C11097 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00108f
C11098 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__inv_1_37/Y 0.00108f
C11099 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.81e-19
C11100 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 2.51e-19
C11101 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_32/HI 0.00508f
C11102 sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__inv_1_27/Y 6.24e-20
C11103 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_48/A 0.0316f
C11104 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_24/A 0.0249f
C11105 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__conb_1_42/HI 9.9e-20
C11106 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# sky130_fd_sc_hd__conb_1_10/HI 4.8e-19
C11107 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q -2.62e-20
C11108 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 1.8e-20
C11109 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0323f
C11110 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 3.23e-21
C11111 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00329f
C11112 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__conb_1_16/HI 8.83e-21
C11113 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__inv_1_50/Y 0.00373f
C11114 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__conb_1_50/HI 0.00699f
C11115 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 4.01e-20
C11116 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# -5.72e-19
C11117 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# -0.0103f
C11118 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__inv_1_33/Y 2.18e-22
C11119 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_51/Y 0.0812f
C11120 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__conb_1_44/HI 4.72e-19
C11121 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_14/Q_N 2.65e-20
C11122 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 8.65e-20
C11123 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# -9.32e-20
C11124 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# 1.38e-20
C11125 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# Reset 3.13e-19
C11126 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.74e-19
C11127 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# -7.17e-20
C11128 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# -1.76e-19
C11129 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0158f
C11130 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# CLOCK_GEN.SR_Op.Q 0.00127f
C11131 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# sky130_fd_sc_hd__inv_1_9/Y 2.73e-20
C11132 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 0.061f
C11133 V_SENSE sky130_fd_sc_hd__inv_1_57/Y 6.82e-19
C11134 sky130_fd_sc_hd__conb_1_10/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 6.65e-20
C11135 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 8.63e-20
C11136 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00186f
C11137 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.31e-19
C11138 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_8/A 0.114f
C11139 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# 2.65e-20
C11140 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 5.05e-19
C11141 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# -6.8e-19
C11142 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.0166f
C11143 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.75e-21
C11144 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 3.54e-21
C11145 sky130_fd_sc_hd__dfbbn_1_2/Q_N FULL_COUNTER.COUNT_SUB_DFF4.Q 1.37e-19
C11146 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -0.00137f
C11147 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0134f
C11148 transmission_gate_9/GN FULL_COUNTER.COUNT_SUB_DFF1.Q 0.141f
C11149 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/Q_N -1.42e-32
C11150 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 2.16e-21
C11151 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 9.14e-20
C11152 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.0595f
C11153 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_1_36/Y 1.07e-21
C11154 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -2.01e-20
C11155 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# -2.18e-19
C11156 sky130_fd_sc_hd__dfbbn_1_48/Q_N V_LOW 1.99e-19
C11157 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_69/Y 2.08e-19
C11158 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q -5.45e-20
C11159 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.917f
C11160 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__inv_1_10/Y 0.0365f
C11161 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.67e-20
C11162 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_67/A 4.24e-20
C11163 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_581_47# -7.91e-19
C11164 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0579f
C11165 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# V_LOW 4.8e-20
C11166 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 5.77e-20
C11167 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_193_47# -0.0319f
C11168 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00245f
C11169 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# V_LOW 2.26e-20
C11170 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q -5.45e-20
C11171 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_1_46/A 0.166f
C11172 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.0165f
C11173 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# sky130_fd_sc_hd__conb_1_5/HI 5.48e-20
C11174 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# 1.11e-20
C11175 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_1_40/Y 1.55e-21
C11176 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_26/HI 5.68e-20
C11177 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_22/Y 0.0932f
C11178 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__conb_1_14/HI 2.33e-20
C11179 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_21/LO 0.00432f
C11180 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -1.61e-19
C11181 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_473_413# -0.00834f
C11182 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# -1.63e-19
C11183 FULL_COUNTER.COUNT_SUB_DFF7.Q V_LOW 2.08f
C11184 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# V_LOW 3.56e-20
C11185 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_1_63/Y 6.08e-22
C11186 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 7.9e-19
C11187 sky130_fd_sc_hd__dfbbn_1_43/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00255f
C11188 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0416f
C11189 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_32/HI 0.0045f
C11190 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_7/HI 2.86e-19
C11191 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 9.31e-20
C11192 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.25e-19
C11193 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__conb_1_19/HI 7.58e-21
C11194 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 2.64e-20
C11195 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_44/A 0.0409f
C11196 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00268f
C11197 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__inv_1_37/Y 9.61e-20
C11198 RISING_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 8.03e-21
C11199 FALLING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 2.14f
C11200 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_1_46/A 0.0662f
C11201 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# 0.00138f
C11202 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 0.131f
C11203 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# sky130_fd_sc_hd__conb_1_32/HI 2e-19
C11204 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# V_LOW 2.26e-20
C11205 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 4.99e-19
C11206 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 9.54e-19
C11207 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 0.00108f
C11208 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# -2.53e-20
C11209 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__conb_1_25/HI 3.27e-21
C11210 sky130_fd_sc_hd__dfbbn_1_30/Q_N RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00112f
C11211 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 8.25e-20
C11212 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00173f
C11213 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__conb_1_35/HI 1.21e-21
C11214 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_891_329# 9.74e-19
C11215 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__conb_1_29/HI 9.82e-19
C11216 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_15/HI 5.95e-20
C11217 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# sky130_fd_sc_hd__inv_1_50/Y 1.07e-21
C11218 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00181f
C11219 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# -6.8e-19
C11220 sky130_fd_sc_hd__inv_8_0/Y Reset 2.36e-19
C11221 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.86e-19
C11222 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0364f
C11223 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# V_LOW 0.0254f
C11224 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 3.39e-19
C11225 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 0.0149f
C11226 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/Q_N -4.24e-20
C11227 sky130_fd_sc_hd__dfbbn_1_18/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0231f
C11228 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 7.4e-19
C11229 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# V_LOW -0.108f
C11230 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# CLOCK_GEN.SR_Op.Q 2.57e-19
C11231 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 9.33e-19
C11232 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.08e-19
C11233 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 7e-19
C11234 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# 2.64e-19
C11235 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.41e-19
C11236 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 2.21e-19
C11237 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_33/Y 2.51e-19
C11238 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 1.38e-19
C11239 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_64/A 0.104f
C11240 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_64/Y 3e-19
C11241 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nor2_1_0/Y 0.705f
C11242 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_44/A 0.00533f
C11243 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.0267f
C11244 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.5e-20
C11245 sky130_fd_sc_hd__conb_1_0/HI V_LOW 0.542f
C11246 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__inv_16_40/Y 0.0451f
C11247 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.39e-19
C11248 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.59e-19
C11249 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_23/Y 0.0731f
C11250 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# V_LOW 0.015f
C11251 sky130_fd_sc_hd__inv_1_60/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 1.12e-21
C11252 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 1.99e-19
C11253 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__conb_1_33/HI -0.0018f
C11254 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_12/HI 0.00923f
C11255 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# 1.11e-20
C11256 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# 1.1e-20
C11257 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# sky130_fd_sc_hd__inv_16_40/Y 0.00501f
C11258 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0119f
C11259 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 7.09e-19
C11260 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0428f
C11261 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 0.0222f
C11262 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# -0.00502f
C11263 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# -0.00242f
C11264 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_12/HI 0.557f
C11265 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__conb_1_31/HI 0.0287f
C11266 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_69/Y 0.059f
C11267 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 8e-21
C11268 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 3.67e-21
C11269 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.00146f
C11270 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_40/Y 1.25e-19
C11271 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00113f
C11272 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# V_LOW 0.00572f
C11273 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 2.89e-19
C11274 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 0.00103f
C11275 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__inv_1_22/Y 5.17e-19
C11276 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_21/LO 0.00758f
C11277 sky130_fd_sc_hd__inv_16_47/Y CLOCK_GEN.SR_Op.Q 0.0295f
C11278 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__conb_1_5/HI 9.5e-20
C11279 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__conb_1_28/HI 2.62e-19
C11280 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# -2.57e-20
C11281 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00586f
C11282 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_67/A 0.0333f
C11283 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.33e-19
C11284 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 0.114f
C11285 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_1_35/Y 8.55e-19
C11286 sky130_fd_sc_hd__inv_16_4/Y V_LOW 0.396f
C11287 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0305f
C11288 sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_16_26/Y 2.23e-21
C11289 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_3/Y 6.34e-20
C11290 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# sky130_fd_sc_hd__conb_1_32/HI 5.07e-19
C11291 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_64/A 0.00389f
C11292 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_46/A 5.3e-20
C11293 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 6.33e-20
C11294 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00122f
C11295 sky130_fd_sc_hd__inv_1_33/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.278f
C11296 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_26/LO 4.68e-21
C11297 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.1e-20
C11298 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# sky130_fd_sc_hd__inv_1_44/A 4.97e-19
C11299 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_29/Y 0.0175f
C11300 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_38/LO 2.03e-19
C11301 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# -0.137f
C11302 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_10/a_381_47# 0.00949f
C11303 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_891_329# 2.92e-19
C11304 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 1.16e-19
C11305 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 5.41e-21
C11306 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# -1.44e-20
C11307 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 0.00363f
C11308 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.0141f
C11309 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.00221f
C11310 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_59/Y 3.08e-20
C11311 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__conb_1_27/HI 1.35e-19
C11312 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_16_41/Y 0.143f
C11313 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_8_1/a_27_47# 0.00239f
C11314 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__conb_1_8/LO 6.67e-21
C11315 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_3/Y 0.0259f
C11316 sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0028f
C11317 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__conb_1_0/HI 2.52e-19
C11318 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# V_LOW 4.8e-20
C11319 sky130_fd_sc_hd__conb_1_36/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 3.39e-19
C11320 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__conb_1_45/HI 0.00245f
C11321 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 8.3e-19
C11322 sky130_fd_sc_hd__conb_1_28/LO FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.88e-20
C11323 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# V_LOW 0.0056f
C11324 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_47/Y 2.37e-20
C11325 sky130_fd_sc_hd__inv_1_47/Y Reset 0.0125f
C11326 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 0.00107f
C11327 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00119f
C11328 FALLING_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 0.82f
C11329 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# V_LOW -2.68e-19
C11330 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 1.72e-19
C11331 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.21e-21
C11332 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0024f
C11333 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 3.57e-20
C11334 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00124f
C11335 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.257f
C11336 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0484f
C11337 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__inv_1_64/Y 6.3e-21
C11338 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.032f
C11339 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_6/HI 1.73e-19
C11340 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# V_LOW 1.38e-19
C11341 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# -6.43e-20
C11342 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# -3.06e-20
C11343 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 5.02e-20
C11344 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# sky130_fd_sc_hd__conb_1_33/HI -0.00248f
C11345 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__conb_1_12/HI 0.0124f
C11346 sky130_fd_sc_hd__inv_1_53/Y CLOCK_GEN.SR_Op.Q 0.00166f
C11347 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 7.69e-20
C11348 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/Q_N -4.33e-20
C11349 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# sky130_fd_sc_hd__conb_1_31/HI 9.52e-19
C11350 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0745f
C11351 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__nand3_1_1/Y 2.22e-20
C11352 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00188f
C11353 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.88e-19
C11354 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_53/A 0.0298f
C11355 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 1.97e-19
C11356 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_67/A 0.00189f
C11357 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00107f
C11358 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_381_47# -2.53e-20
C11359 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# 0.00122f
C11360 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__conb_1_24/HI 5.87e-20
C11361 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__conb_1_28/HI -6.57e-19
C11362 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__conb_1_5/HI 4.88e-20
C11363 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.024f
C11364 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0174f
C11365 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.67e-21
C11366 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 8e-21
C11367 sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__inv_1_31/Y 9.11e-20
C11368 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_56/Y 2.84e-19
C11369 sky130_fd_sc_hd__conb_1_50/LO V_LOW 0.0522f
C11370 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00408f
C11371 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.38e-19
C11372 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__inv_1_35/Y 0.0137f
C11373 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_29/A 0.0188f
C11374 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_7/LO 0.00511f
C11375 sky130_fd_sc_hd__inv_1_60/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00454f
C11376 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__conb_1_2/HI 3.95e-19
C11377 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_41/HI 0.0251f
C11378 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 0.0296f
C11379 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.00808f
C11380 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 8.95e-21
C11381 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__inv_1_44/A 0.00388f
C11382 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# sky130_fd_sc_hd__conb_1_20/HI 3.89e-19
C11383 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# V_LOW 0.00883f
C11384 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# Reset 0.00243f
C11385 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00257f
C11386 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1_19/HI 0.00808f
C11387 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_381_47# 0.00465f
C11388 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_1/Y 0.024f
C11389 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.4e-19
C11390 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00222f
C11391 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# -0.00524f
C11392 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_891_329# -0.00159f
C11393 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 3.44e-19
C11394 sky130_fd_sc_hd__conb_1_10/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0262f
C11395 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 7.69e-19
C11396 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__dfbbn_1_27/Q_N 5.89e-19
C11397 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__inv_1_60/Y 0.0309f
C11398 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 3.45e-19
C11399 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0844f
C11400 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand3_1_2/Y 1.38e-21
C11401 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_1_14/Y 8.46e-19
C11402 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# sky130_fd_sc_hd__conb_1_0/HI 2.43e-19
C11403 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0152f
C11404 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__inv_1_31/Y 3.94e-20
C11405 sky130_fd_sc_hd__inv_1_5/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 8.43e-19
C11406 sky130_fd_sc_hd__dfbbn_1_49/a_581_47# sky130_fd_sc_hd__conb_1_45/HI 0.00213f
C11407 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.0152f
C11408 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 0.00964f
C11409 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_16_2/Y 0.0132f
C11410 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# 2.46e-19
C11411 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00251f
C11412 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00135f
C11413 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_19/HI 2.01e-21
C11414 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__conb_1_11/HI 1.76e-20
C11415 FALLING_COUNTER.COUNT_SUB_DFF10.Q V_LOW 2.94f
C11416 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 4.36e-19
C11417 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00635f
C11418 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_29/HI 1.13e-22
C11419 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# sky130_fd_sc_hd__inv_1_10/Y 1.04e-19
C11420 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__conb_1_50/HI 7.69e-19
C11421 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.016f
C11422 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__conb_1_6/HI -7.08e-20
C11423 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.54e-22
C11424 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0.00123f
C11425 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 1.39e-19
C11426 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 0.00206f
C11427 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_43/Q_N 4.52e-21
C11428 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# 6.95e-21
C11429 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_53/Y 4.81e-21
C11430 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_1_28/Y 0.00373f
C11431 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.13e-21
C11432 sky130_fd_sc_hd__dfbbn_1_4/Q_N FULL_COUNTER.COUNT_SUB_DFF7.Q 0.033f
C11433 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__conb_1_48/LO 0.0037f
C11434 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__conb_1_7/HI 1.44e-21
C11435 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/Q_N -9.56e-20
C11436 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_2_0/A 0.0161f
C11437 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_46/A 0.498f
C11438 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# sky130_fd_sc_hd__inv_1_41/Y 3.39e-19
C11439 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_1_21/Y 0.00421f
C11440 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 9.25e-20
C11441 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# -6.43e-20
C11442 sky130_fd_sc_hd__nand2_8_9/A FULL_COUNTER.COUNT_SUB_DFF2.Q 2.21e-19
C11443 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# -0.0147f
C11444 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 2.39e-21
C11445 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.46e-19
C11446 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# -1.44e-20
C11447 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0151f
C11448 sky130_fd_sc_hd__inv_1_40/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 2.71e-21
C11449 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_193_47# -0.236f
C11450 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 3.01e-21
C11451 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 4.13e-19
C11452 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_25/Y 1.77e-20
C11453 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 2e-19
C11454 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_21/Y 0.0016f
C11455 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__inv_16_41/Y 0.136f
C11456 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 7.48e-21
C11457 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 6.82e-20
C11458 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_7/LO 4.17e-19
C11459 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__conb_1_23/LO 9.17e-19
C11460 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 1.67e-21
C11461 FALLING_COUNTER.COUNT_SUB_DFF13.Q V_LOW 1.55f
C11462 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# V_LOW 3.56e-20
C11463 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__conb_1_32/HI 1.58e-20
C11464 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# 3.53e-19
C11465 sky130_fd_sc_hd__inv_1_65/A FULL_COUNTER.COUNT_SUB_DFF1.Q 5.78e-20
C11466 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 7.23e-21
C11467 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 3.07e-19
C11468 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.39e-19
C11469 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__nand2_8_4/Y 0.0169f
C11470 sky130_fd_sc_hd__nand2_8_4/a_27_47# Reset 0.0468f
C11471 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# Reset 1.7e-19
C11472 transmission_gate_9/GN FULL_COUNTER.COUNT_SUB_DFF0.Q 0.143f
C11473 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_44/A 5.39e-20
C11474 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# CLOCK_GEN.SR_Op.Q 0.034f
C11475 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# V_LOW 1.38e-19
C11476 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 9.57e-20
C11477 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 3.85e-20
C11478 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00483f
C11479 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0163f
C11480 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_19/Y 4.56e-19
C11481 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.21e-19
C11482 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# -0.00385f
C11483 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_4/HI 0.0301f
C11484 sky130_fd_sc_hd__conb_1_48/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00407f
C11485 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_891_329# -2.2e-20
C11486 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# -0.00859f
C11487 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 5.49e-20
C11488 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00697f
C11489 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__inv_1_39/Y 0.0671f
C11490 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# V_LOW 2.26e-20
C11491 sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__conb_1_0/HI 4.38e-20
C11492 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_40/HI 0.494f
C11493 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0128f
C11494 sky130_fd_sc_hd__inv_16_6/Y V_LOW 0.295f
C11495 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__inv_1_8/Y 1.83e-19
C11496 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0652f
C11497 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__inv_16_40/Y 0.0023f
C11498 sky130_fd_sc_hd__dfbbn_1_41/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0152f
C11499 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__inv_1_61/Y 6.69e-20
C11500 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__conb_1_4/HI 0.0036f
C11501 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0225f
C11502 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__inv_1_38/Y 6.65e-20
C11503 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_29/HI 0.00556f
C11504 sky130_fd_sc_hd__dfbbn_1_26/a_581_47# sky130_fd_sc_hd__conb_1_50/HI 1.14e-19
C11505 sky130_fd_sc_hd__nand2_1_1/a_113_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.61e-19
C11506 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 2.38e-19
C11507 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_557_413# -3.67e-20
C11508 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# -6.29e-19
C11509 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_16/LO 2.73e-19
C11510 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_1_39/Y 0.00143f
C11511 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.49e-21
C11512 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_24/A 0.0102f
C11513 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0911f
C11514 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_16_41/Y 0.571f
C11515 RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0083f
C11516 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# sky130_fd_sc_hd__conb_1_47/HI 8.33e-19
C11517 sky130_fd_sc_hd__conb_1_38/LO FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00218f
C11518 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00102f
C11519 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# sky130_fd_sc_hd__inv_1_28/Y 5.83e-21
C11520 sky130_fd_sc_hd__inv_16_40/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0335f
C11521 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 3.8e-21
C11522 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 4.48e-19
C11523 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 0.0236f
C11524 sky130_fd_sc_hd__inv_16_33/Y V_LOW 0.176f
C11525 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_15/LO 0.00178f
C11526 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# -0.11f
C11527 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_64/A 0.0234f
C11528 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__inv_1_21/Y 1.74e-20
C11529 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__inv_1_39/Y 0.0117f
C11530 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__inv_1_44/A 0.0067f
C11531 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0396f
C11532 RISING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00404f
C11533 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_16_40/Y 0.587f
C11534 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__conb_1_15/HI 7.44e-20
C11535 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# sky130_fd_sc_hd__conb_1_10/HI 2.66e-20
C11536 FALLING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 1.34e-20
C11537 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_26/Y 1.63e-20
C11538 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00302f
C11539 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.119f
C11540 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0943f
C11541 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__inv_1_60/Y 2.21e-20
C11542 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# sky130_fd_sc_hd__inv_1_55/Y 0.00202f
C11543 sky130_fd_sc_hd__inv_16_6/Y sky130_fd_sc_hd__inv_16_9/Y 0.00249f
C11544 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 5.12e-21
C11545 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_23/HI 0.427f
C11546 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_15/HI -0.0788f
C11547 V_HIGH FULL_COUNTER.COUNT_SUB_DFF7.Q 0.919f
C11548 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__inv_1_43/Y 1.32e-20
C11549 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__conb_1_8/HI -0.00252f
C11550 sky130_fd_sc_hd__inv_16_52/A sky130_fd_sc_hd__inv_16_50/A 0.00257f
C11551 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_48/A 0.722f
C11552 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# -0.00155f
C11553 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# -0.0152f
C11554 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 6.71e-19
C11555 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 4.56e-21
C11556 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_16_2/Y 0.00595f
C11557 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# V_LOW 0.0093f
C11558 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# V_LOW -0.00121f
C11559 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_34/HI 5.47e-20
C11560 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_891_329# -2.2e-20
C11561 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# -0.00853f
C11562 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# CLOCK_GEN.SR_Op.Q 7.69e-20
C11563 sky130_fd_sc_hd__inv_1_60/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.69e-19
C11564 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_29/Y 8.63e-19
C11565 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# V_LOW 0.019f
C11566 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# V_LOW 0.006f
C11567 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# V_LOW -0.00121f
C11568 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__inv_1_30/Y 6.82e-20
C11569 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__dfbbn_1_27/a_381_47# 1.74e-19
C11570 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__conb_1_7/HI 0.00937f
C11571 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.08e-19
C11572 FULL_COUNTER.COUNT_SUB_DFF18.Q sky130_fd_sc_hd__conb_1_11/HI 0.00382f
C11573 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# -0.00592f
C11574 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# sky130_fd_sc_hd__inv_16_41/Y 5.67e-19
C11575 sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 6.32e-19
C11576 sky130_fd_sc_hd__inv_16_33/Y sky130_fd_sc_hd__inv_16_9/Y 0.0616f
C11577 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# V_LOW -0.0133f
C11578 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 0.00638f
C11579 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# V_LOW -0.00266f
C11580 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_15/HI 9.92e-21
C11581 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__conb_1_39/HI 1.63e-20
C11582 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# sky130_fd_sc_hd__inv_1_8/Y 5.8e-19
C11583 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0646f
C11584 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_16_19/Y 2.39e-19
C11585 FALLING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 3.93f
C11586 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_42/Y 0.00807f
C11587 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 2.47e-20
C11588 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__inv_1_38/Y 2e-19
C11589 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 1.37e-19
C11590 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_29/HI 0.0185f
C11591 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# V_LOW 0.0358f
C11592 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_1_32/Y 5.2e-20
C11593 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_50/HI 6.13e-20
C11594 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__conb_1_26/HI 4.32e-20
C11595 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# V_LOW 0.00471f
C11596 sky130_fd_sc_hd__inv_1_62/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.237f
C11597 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_49/Y 1.45f
C11598 sky130_fd_sc_hd__conb_1_0/HI V_HIGH 5.97e-19
C11599 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.14e-19
C11600 sky130_fd_sc_hd__inv_2_0/A FULL_COUNTER.COUNT_SUB_DFF2.Q 0.124f
C11601 FULL_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.52e-19
C11602 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 7.16e-19
C11603 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_28/LO 5.25e-20
C11604 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_23/A 1.42e-19
C11605 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__conb_1_51/HI 0.0024f
C11606 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 7.51e-21
C11607 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI 0.02f
C11608 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_55/A 0.614f
C11609 sky130_fd_sc_hd__nand2_8_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.22e-19
C11610 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# sky130_fd_sc_hd__inv_1_44/A 2.96e-19
C11611 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_64/Y 0.00133f
C11612 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_3/A 0.0141f
C11613 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0482f
C11614 sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.14f
C11615 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.332f
C11616 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# V_LOW -9.15e-19
C11617 sky130_fd_sc_hd__conb_1_30/HI V_LOW 0.185f
C11618 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__inv_1_14/Y 1.6e-19
C11619 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# sky130_fd_sc_hd__inv_16_42/Y 6.65e-21
C11620 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 2.13e-20
C11621 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# sky130_fd_sc_hd__conb_1_6/HI 0.00369f
C11622 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_5/Y 0.123f
C11623 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_14/Y 0.0749f
C11624 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.027f
C11625 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0453f
C11626 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00438f
C11627 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00871f
C11628 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.62e-21
C11629 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 4.62e-19
C11630 sky130_fd_sc_hd__inv_1_55/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.138f
C11631 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_49/Y 0.368f
C11632 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 1.25e-20
C11633 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_33/HI 4.84e-20
C11634 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/Q_N 9.65e-21
C11635 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 7.38e-22
C11636 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_8_8/A 0.00868f
C11637 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 0.00851f
C11638 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.37e-20
C11639 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 5.18e-19
C11640 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -0.0037f
C11641 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# -0.012f
C11642 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 0.00124f
C11643 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__conb_1_50/HI 0.012f
C11644 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_941_21# 2.39e-19
C11645 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_67/A 0.014f
C11646 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 4.31e-19
C11647 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__conb_1_17/HI 0.002f
C11648 sky130_fd_sc_hd__dfbbn_1_35/Q_N CLOCK_GEN.SR_Op.Q 0.0215f
C11649 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# -0.00592f
C11650 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 7.86e-21
C11651 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# V_LOW -6.55e-19
C11652 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__inv_1_64/A 0.00586f
C11653 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_32/Y 0.0889f
C11654 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# V_LOW -1.39e-35
C11655 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 3.55e-19
C11656 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.8e-20
C11657 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_647_21# -1.69e-19
C11658 V_SENSE sky130_fd_sc_hd__fill_4_194/VPB 0.0211f
C11659 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 9.58e-21
C11660 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# V_LOW 4.8e-20
C11661 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_891_329# 0.00143f
C11662 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# V_LOW -0.00795f
C11663 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__conb_1_37/HI 5.87e-21
C11664 sky130_fd_sc_hd__conb_1_5/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 1.05e-20
C11665 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0354f
C11666 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0219f
C11667 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 5.54e-19
C11668 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__conb_1_24/HI 0.0278f
C11669 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0127f
C11670 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__inv_1_13/Y 2.46e-22
C11671 sky130_fd_sc_hd__conb_1_45/HI sky130_fd_sc_hd__inv_1_61/Y 0.133f
C11672 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_66/Y 6.91e-19
C11673 sky130_fd_sc_hd__inv_1_35/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 5.99e-21
C11674 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0282f
C11675 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0248f
C11676 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# -0.012f
C11677 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -0.0133f
C11678 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__conb_1_38/HI 4.64e-19
C11679 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 4.11e-19
C11680 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# V_LOW -6.55e-19
C11681 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 6.1e-19
C11682 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_51/A 0.111f
C11683 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 0.0079f
C11684 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0198f
C11685 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.123f
C11686 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_24/HI 1.63e-19
C11687 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__conb_1_44/HI 0.00118f
C11688 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__conb_1_48/HI 0.00983f
C11689 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00638f
C11690 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_46/A 0.00133f
C11691 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# V_LOW -0.00371f
C11692 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0421f
C11693 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0016f
C11694 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.03e-20
C11695 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00163f
C11696 sky130_fd_sc_hd__conb_1_13/HI V_LOW 0.148f
C11697 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 2.73e-20
C11698 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__nand2_8_9/A 9.55e-19
C11699 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__inv_1_14/Y 3.29e-19
C11700 V_SENSE sky130_fd_sc_hd__conb_1_49/HI 0.00142f
C11701 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 0.00353f
C11702 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__inv_1_33/Y 0.0376f
C11703 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 0.014f
C11704 sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF12.Q 0.125f
C11705 sky130_fd_sc_hd__conb_1_38/HI V_LOW 0.178f
C11706 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 6.17e-20
C11707 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 6.17e-20
C11708 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 1.74e-19
C11709 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 1.74e-19
C11710 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__conb_1_24/LO 0.0015f
C11711 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 1.6e-19
C11712 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.0023f
C11713 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 8.08e-19
C11714 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_0/Y 0.408f
C11715 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0202f
C11716 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__conb_1_0/HI 2.45e-20
C11717 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# V_LOW -0.109f
C11718 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00333f
C11719 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# -0.00591f
C11720 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# -6.43e-20
C11721 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__nor2_1_0/Y 2.44e-21
C11722 sky130_fd_sc_hd__nand3_1_0/Y CLOCK_GEN.SR_Op.Q 0.0908f
C11723 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# -2.57e-20
C11724 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 9.17e-22
C11725 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 2.68e-20
C11726 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 1.15e-22
C11727 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__conb_1_50/HI 0.00232f
C11728 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_35/HI 0.0177f
C11729 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__conb_1_40/HI 2.07e-19
C11730 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 4.12e-19
C11731 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__conb_1_17/HI 9.55e-19
C11732 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/Q_N -6.48e-19
C11733 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.22e-21
C11734 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 8.51e-20
C11735 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF12.Q -2.62e-20
C11736 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# V_LOW 0.022f
C11737 sky130_fd_sc_hd__dfbbn_1_10/Q_N V_LOW -0.00103f
C11738 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 2.93e-20
C11739 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 6.21e-20
C11740 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_941_21# -3.07e-19
C11741 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# -2.37e-19
C11742 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 3.71e-19
C11743 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_581_47# -7.91e-19
C11744 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 0.0155f
C11745 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 4.51e-22
C11746 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_20/HI 0.00112f
C11747 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 8.77e-19
C11748 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 0.0126f
C11749 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 1.45e-19
C11750 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 6.87e-20
C11751 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 1.45e-19
C11752 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 6.87e-20
C11753 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00288f
C11754 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00819f
C11755 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0619f
C11756 V_SENSE sky130_fd_sc_hd__fill_4_184/VPB 0.0211f
C11757 sky130_fd_sc_hd__conb_1_51/HI CLOCK_GEN.SR_Op.Q 6.37e-19
C11758 RISING_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF6.Q 1.71f
C11759 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 9.4e-19
C11760 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_26/Y 0.0117f
C11761 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 1.87e-19
C11762 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 8.29e-20
C11763 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__conb_1_24/HI 0.00254f
C11764 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_52/A 0.0192f
C11765 sky130_fd_sc_hd__inv_1_39/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 5.74e-22
C11766 sky130_fd_sc_hd__conb_1_39/HI V_LOW 0.176f
C11767 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_16_40/Y 5.72e-20
C11768 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_64/Y 1.57e-19
C11769 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 9.2e-19
C11770 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.0026f
C11771 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 6e-20
C11772 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# V_LOW 0.00247f
C11773 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# sky130_fd_sc_hd__conb_1_50/HI 1.2e-19
C11774 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0343f
C11775 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__conb_1_9/HI 0.00281f
C11776 sky130_fd_sc_hd__dfbbn_1_3/a_581_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00101f
C11777 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# -9.41e-19
C11778 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 0.00122f
C11779 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_557_413# -3.67e-20
C11780 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# -0.00717f
C11781 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_891_329# -2.46e-19
C11782 sky130_fd_sc_hd__inv_1_65/A FULL_COUNTER.COUNT_SUB_DFF0.Q 1.28e-20
C11783 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0414f
C11784 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.85e-20
C11785 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_8_0/Y 0.0295f
C11786 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 4.01e-19
C11787 sky130_fd_sc_hd__dfbbn_1_16/Q_N V_LOW -0.00452f
C11788 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_20/A 5.07e-19
C11789 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 9.06e-20
C11790 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_24/A 7.15e-21
C11791 sky130_fd_sc_hd__inv_1_45/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.107f
C11792 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_13/LO 0.0144f
C11793 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0162f
C11794 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00111f
C11795 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0452f
C11796 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_14/HI 0.0307f
C11797 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__conb_1_10/HI 7.44e-20
C11798 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__conb_1_48/HI -1.93e-19
C11799 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0402f
C11800 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__conb_1_39/HI 0.00166f
C11801 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0.0573f
C11802 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_1_5/Y 1.01e-19
C11803 sky130_fd_sc_hd__inv_16_6/A RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0297f
C11804 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__inv_1_50/Y 0.0143f
C11805 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_46/A 9.76e-22
C11806 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# -0.00161f
C11807 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 0.00177f
C11808 sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 8.14e-21
C11809 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 4.83e-19
C11810 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# 8.44e-19
C11811 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__inv_1_27/Y 1.32e-21
C11812 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0267f
C11813 RISING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0016f
C11814 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 0.0365f
C11815 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_381_47# -3.79e-20
C11816 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# -4.66e-20
C11817 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.03e-20
C11818 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# sky130_fd_sc_hd__inv_1_0/Y 5.77e-20
C11819 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 6.55e-20
C11820 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 0.0353f
C11821 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# V_LOW -9.94e-19
C11822 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_46/A 0.0113f
C11823 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__inv_16_40/Y 0.0186f
C11824 sky130_fd_sc_hd__conb_1_3/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 8.23e-19
C11825 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_25/LO 1.3e-20
C11826 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__inv_1_41/Y 0.00918f
C11827 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00372f
C11828 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_1_59/Y 0.317f
C11829 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 3.16e-21
C11830 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 2.51e-22
C11831 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__conb_1_35/HI 0.00252f
C11832 FULL_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0355f
C11833 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__conb_1_40/HI -0.00656f
C11834 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.75e-21
C11835 RISING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.09f
C11836 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.014f
C11837 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0379f
C11838 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# V_LOW 3.56e-20
C11839 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.07e-19
C11840 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__conb_1_8/HI 3.34e-21
C11841 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# -9.52e-20
C11842 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_1_49/Y 0.0465f
C11843 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# V_LOW 0.0102f
C11844 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 0.00491f
C11845 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# -7.17e-20
C11846 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# -1.66e-19
C11847 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 2.1e-19
C11848 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 0.00196f
C11849 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 4.99e-19
C11850 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 9.54e-19
C11851 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0.00108f
C11852 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_5/A 0.0488f
C11853 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__conb_1_26/HI 1.61e-19
C11854 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00113f
C11855 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0047f
C11856 RISING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 1.63f
C11857 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_51/HI 0.02f
C11858 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 3.1e-20
C11859 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# 5.14e-19
C11860 sky130_fd_sc_hd__inv_1_35/Y sky130_fd_sc_hd__inv_16_41/Y 0.0249f
C11861 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.35e-19
C11862 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# sky130_fd_sc_hd__inv_1_26/Y 0.00152f
C11863 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0882f
C11864 sky130_fd_sc_hd__dfbbn_1_5/Q_N FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0256f
C11865 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 2.55e-19
C11866 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.0399f
C11867 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__conb_1_27/HI 8.12e-22
C11868 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__inv_1_2/Y 1.07e-20
C11869 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# V_LOW 0.0233f
C11870 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_30/Y 9.48e-21
C11871 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.76e-20
C11872 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.63e-20
C11873 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# -0.00497f
C11874 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_1_30/Y 1.39e-19
C11875 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00588f
C11876 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_7/HI 0.00341f
C11877 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00293f
C11878 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 3.81e-20
C11879 V_SENSE sky130_fd_sc_hd__inv_16_9/A 0.17f
C11880 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__conb_1_3/HI -0.00164f
C11881 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__nand3_1_2/Y 5.97e-19
C11882 sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00146f
C11883 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.07e-19
C11884 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# V_LOW 0.0292f
C11885 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__inv_1_9/Y 0.122f
C11886 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_1_33/Y 0.0014f
C11887 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__conb_1_0/HI 0.00624f
C11888 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 3.89e-19
C11889 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 2.45e-20
C11890 sky130_fd_sc_hd__nor2_1_0/Y Reset 0.0843f
C11891 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 6.25e-21
C11892 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.2e-19
C11893 sky130_fd_sc_hd__conb_1_47/LO V_LOW 0.0857f
C11894 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_2_0/A 0.0459f
C11895 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__inv_16_42/Y 0.051f
C11896 sky130_fd_sc_hd__conb_1_34/HI V_LOW 0.131f
C11897 FULL_COUNTER.COUNT_SUB_DFF2.Q V_LOW 0.814f
C11898 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__conb_1_14/HI -0.0119f
C11899 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 1.01e-19
C11900 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_9/HI 6.05e-19
C11901 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.27e-19
C11902 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__inv_1_63/Y 0.0209f
C11903 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00493f
C11904 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 0.034f
C11905 V_SENSE sky130_fd_sc_hd__inv_16_22/A 0.156f
C11906 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# 3.94e-21
C11907 sky130_fd_sc_hd__conb_1_25/LO V_LOW 0.0513f
C11908 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0452f
C11909 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/Q_N 0.00144f
C11910 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_24/A 0.0308f
C11911 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# Reset 0.00429f
C11912 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_23/HI 0.0142f
C11913 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# 0.0248f
C11914 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 3.42e-19
C11915 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.08e-20
C11916 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.011f
C11917 sky130_fd_sc_hd__conb_1_36/LO V_LOW 0.0934f
C11918 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__conb_1_31/HI 0.00475f
C11919 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__conb_1_2/HI 0.0106f
C11920 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__inv_1_41/Y 0.00129f
C11921 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_34/HI 0.264f
C11922 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00463f
C11923 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 2.32e-20
C11924 sky130_fd_sc_hd__conb_1_9/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 0.016f
C11925 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.83e-20
C11926 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00147f
C11927 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0438f
C11928 sky130_fd_sc_hd__conb_1_14/LO V_LOW 0.0604f
C11929 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_891_329# 9.74e-19
C11930 sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_16_23/Y 0.161f
C11931 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_64/A 1.42e-21
C11932 Reset sky130_fd_sc_hd__inv_1_64/A 0.0112f
C11933 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# -0.00336f
C11934 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# -3.79e-20
C11935 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__inv_1_1/Y 4.3e-21
C11936 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_581_47# -2.6e-20
C11937 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 3.5e-20
C11938 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00854f
C11939 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# 0.00185f
C11940 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00511f
C11941 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__inv_1_40/Y 0.00103f
C11942 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 1.16e-19
C11943 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.69e-19
C11944 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_45/HI 0.0129f
C11945 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_557_413# -3.67e-20
C11946 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_891_329# -2.46e-19
C11947 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# -0.0234f
C11948 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__conb_1_38/HI 8.37e-20
C11949 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__inv_2_0/A 3.63e-20
C11950 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_45/Y 0.00346f
C11951 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_40/a_193_47# 3.23e-19
C11952 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.37e-20
C11953 sky130_fd_sc_hd__inv_16_15/Y V_LOW 0.306f
C11954 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.00449f
C11955 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 3.85e-19
C11956 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 7.76e-19
C11957 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 9.18e-20
C11958 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_32/HI 1.81e-20
C11959 sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00497f
C11960 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# V_LOW 0.00358f
C11961 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 0.0115f
C11962 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_16_4/Y 0.0919f
C11963 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.0184f
C11964 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# V_LOW 0.00498f
C11965 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# -0.00141f
C11966 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# -0.00367f
C11967 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -9.88e-20
C11968 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# -6.23e-21
C11969 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__inv_1_30/Y 2.74e-19
C11970 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.67e-20
C11971 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.26e-21
C11972 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/Q_N 7.66e-19
C11973 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__inv_1_60/Y 0.00848f
C11974 sky130_fd_sc_hd__conb_1_2/HI V_LOW 0.152f
C11975 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_381_47# -2.53e-20
C11976 sky130_fd_sc_hd__inv_16_31/Y sky130_fd_sc_hd__inv_16_7/A 0.0736f
C11977 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# V_LOW 2.94e-20
C11978 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 2.32e-20
C11979 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__inv_16_40/Y 0.00226f
C11980 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__inv_16_42/Y 0.0202f
C11981 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0823f
C11982 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 0.0773f
C11983 RISING_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.946f
C11984 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 0.281f
C11985 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 1.33e-19
C11986 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_29/Y 0.00167f
C11987 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# 9.52e-19
C11988 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 4.02e-20
C11989 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 2.99e-20
C11990 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.72e-19
C11991 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_2_0/A 5.91e-20
C11992 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00176f
C11993 V_SENSE sky130_fd_sc_hd__inv_16_51/A 0.431f
C11994 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 8.63e-20
C11995 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 3.92e-20
C11996 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__inv_1_9/Y 0.00314f
C11997 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_46/A 0.148f
C11998 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_1_43/Y 0.0031f
C11999 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# sky130_fd_sc_hd__inv_1_27/Y 7.05e-19
C12000 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# Reset 0.0014f
C12001 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# sky130_fd_sc_hd__conb_1_23/HI 3.17e-20
C12002 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_31/HI 9.21e-21
C12003 sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__inv_1_27/Y 4.84e-20
C12004 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# 0.0108f
C12005 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.85e-19
C12006 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_473_413# 0.00533f
C12007 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_28/LO 0.0624f
C12008 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0404f
C12009 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__conb_1_2/HI -1.28e-19
C12010 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_1_41/Y 0.0232f
C12011 sky130_fd_sc_hd__inv_16_41/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.114f
C12012 sky130_fd_sc_hd__inv_1_30/Y sky130_fd_sc_hd__inv_1_29/Y 1.48e-19
C12013 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__inv_1_13/Y 0.00721f
C12014 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_891_329# -2.46e-19
C12015 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# -0.00311f
C12016 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_557_413# -3.67e-20
C12017 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_891_329# -2.2e-20
C12018 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# -0.00788f
C12019 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 4.27e-19
C12020 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__inv_1_32/Y 3.99e-20
C12021 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0287f
C12022 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# V_LOW 0.00864f
C12023 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 2.5e-19
C12024 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0522f
C12025 sky130_fd_sc_hd__conb_1_25/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 1.7e-20
C12026 sky130_fd_sc_hd__conb_1_26/HI V_LOW 0.146f
C12027 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 0.0262f
C12028 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_1_1/Y 8.03e-19
C12029 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 7.69e-19
C12030 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__inv_1_69/Y 4.4e-19
C12031 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.23e-20
C12032 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.72e-19
C12033 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# -5.42e-19
C12034 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00558f
C12035 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 9.21e-20
C12036 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 0.00523f
C12037 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 1.01e-20
C12038 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_381_47# 0.00117f
C12039 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_44/A 0.153f
C12040 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00492f
C12041 sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0823f
C12042 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_33/Y 0.158f
C12043 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__inv_1_50/Y 1.01e-19
C12044 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 1.96e-20
C12045 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 4.34e-19
C12046 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__conb_1_39/LO 1.64e-20
C12047 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__inv_16_41/Y 0.272f
C12048 sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__inv_1_2/Y 5.85e-22
C12049 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# V_LOW 0.00667f
C12050 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__inv_1_36/Y 8.33e-21
C12051 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_891_329# 1.69e-21
C12052 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__conb_1_31/HI 1.34e-21
C12053 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# -3.79e-20
C12054 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# -4.66e-20
C12055 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 3.44e-20
C12056 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand2_8_4/Y 0.0215f
C12057 sky130_fd_sc_hd__nand3_1_2/Y Reset 0.111f
C12058 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__inv_1_32/Y 2.32e-19
C12059 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# V_LOW -0.00121f
C12060 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# V_LOW -0.00266f
C12061 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# V_LOW -2.78e-35
C12062 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0254f
C12063 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_1_59/Y 0.00417f
C12064 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# V_LOW 3.56e-20
C12065 sky130_fd_sc_hd__conb_1_18/LO RISING_COUNTER.COUNT_SUB_DFF15.Q 0.021f
C12066 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -0.00932f
C12067 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# -0.012f
C12068 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__conb_1_28/HI 9.67e-20
C12069 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# Reset 0.0116f
C12070 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__inv_1_44/A 0.0269f
C12071 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_6/HI 0.0115f
C12072 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# 0.0063f
C12073 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 8.76e-23
C12074 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# -1.44e-20
C12075 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 3.39e-19
C12076 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# V_LOW 1.38e-19
C12077 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.28e-19
C12078 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# V_LOW -0.00151f
C12079 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__inv_16_42/Y 0.0294f
C12080 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__nor2_1_0/Y 0.00217f
C12081 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_16_41/Y 2.33e-20
C12082 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5e-19
C12083 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 2.05e-19
C12084 sky130_fd_sc_hd__inv_1_57/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0657f
C12085 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 1.51e-20
C12086 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 8.15e-20
C12087 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 8.15e-20
C12088 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 1.51e-20
C12089 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# 0.00218f
C12090 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 9.14e-19
C12091 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 7.34e-19
C12092 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 1e-19
C12093 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0126f
C12094 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__inv_1_29/Y 1.78e-20
C12095 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.22e-21
C12096 FALLING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 6.05e-20
C12097 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_1_43/Y 4.39e-20
C12098 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 8.68e-19
C12099 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__inv_1_63/Y 0.046f
C12100 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_64/A 0.00106f
C12101 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# 1.22e-20
C12102 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__inv_16_41/Y 1.3e-19
C12103 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_2/LO 1.26e-20
C12104 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_19/A 0.0948f
C12105 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__conb_1_37/HI 6.75e-19
C12106 sky130_fd_sc_hd__inv_1_40/Y RISING_COUNTER.COUNT_SUB_DFF8.Q 0.264f
C12107 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0362f
C12108 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.00169f
C12109 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# -0.0847f
C12110 sky130_fd_sc_hd__dfbbn_1_36/Q_N Reset 2.88e-21
C12111 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# V_LOW 3.56e-20
C12112 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/Q_N 0.0265f
C12113 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 2.69e-20
C12114 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 5.29e-20
C12115 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# 0.00104f
C12116 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.0366f
C12117 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.00609f
C12118 sky130_fd_sc_hd__inv_16_55/Y sky130_fd_sc_hd__inv_16_48/A 0.00169f
C12119 sky130_fd_sc_hd__inv_16_51/Y sky130_fd_sc_hd__inv_16_50/A 0.225f
C12120 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 8.74e-20
C12121 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__conb_1_2/HI -2.17e-19
C12122 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00938f
C12123 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 8.15e-20
C12124 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 2.62e-20
C12125 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 2.78e-19
C12126 sky130_fd_sc_hd__inv_16_27/Y V_LOW 0.14f
C12127 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# -0.00385f
C12128 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__inv_1_32/Y 6.08e-21
C12129 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00994f
C12130 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# V_LOW 6.02e-20
C12131 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# sky130_fd_sc_hd__inv_1_28/Y 0.0015f
C12132 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0161f
C12133 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0272f
C12134 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# V_LOW 0.00546f
C12135 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__inv_1_1/Y 0.00116f
C12136 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.87f
C12137 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 3.47e-19
C12138 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_16_40/Y 0.00121f
C12139 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 0.032f
C12140 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 5.76e-19
C12141 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_61/Y 6.56e-19
C12142 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__inv_1_30/Y 0.00186f
C12143 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# sky130_fd_sc_hd__inv_1_50/Y 5.83e-21
C12144 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_891_329# -2.2e-20
C12145 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# -0.00859f
C12146 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__inv_16_41/Y 0.0402f
C12147 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00353f
C12148 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# sky130_fd_sc_hd__inv_1_36/Y 4.67e-21
C12149 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_1_35/Y 0.0198f
C12150 sky130_fd_sc_hd__dfbbn_1_20/Q_N V_LOW -0.00509f
C12151 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.00687f
C12152 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0283f
C12153 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/Q_N -9.56e-20
C12154 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# V_LOW 0.00466f
C12155 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.37e-20
C12156 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0352f
C12157 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__inv_1_69/Y 8.51e-19
C12158 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_16_40/Y 0.326f
C12159 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# -0.00497f
C12160 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# -2.57e-20
C12161 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_55/Y 0.316f
C12162 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__inv_1_44/A 7.69e-20
C12163 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_26/HI 0.0672f
C12164 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__inv_16_41/Y 0.0322f
C12165 FULL_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.27f
C12166 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# V_LOW 2.94e-20
C12167 V_SENSE sky130_fd_sc_hd__inv_16_19/Y 0.00205f
C12168 sky130_fd_sc_hd__inv_1_22/Y V_LOW 0.132f
C12169 sky130_fd_sc_hd__dfbbn_1_3/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6e-20
C12170 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_891_329# -2.2e-20
C12171 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# -3.48e-20
C12172 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 2.56e-19
C12173 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 2.56e-19
C12174 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_34/HI 0.0278f
C12175 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_0/a_381_47# 6.87e-21
C12176 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_16_50/A 0.0272f
C12177 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.4e-19
C12178 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.672f
C12179 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_1_43/Y 3.48e-21
C12180 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_56/A 0.208f
C12181 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__conb_1_30/LO 2.36e-20
C12182 sky130_fd_sc_hd__inv_1_52/A V_LOW 0.23f
C12183 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 9.32e-19
C12184 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 6.42e-21
C12185 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_55/Y 0.302f
C12186 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00136f
C12187 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00506f
C12188 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_16_4/Y 0.0103f
C12189 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# V_LOW 2.26e-20
C12190 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 9.23e-19
C12191 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00161f
C12192 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_44/A 2.01e-20
C12193 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 9.26e-19
C12194 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_48/A 0.00788f
C12195 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8_9/A 0.00141f
C12196 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.87e-21
C12197 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 6.35e-19
C12198 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_19/Y 0.00146f
C12199 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 1.39e-21
C12200 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# -0.00375f
C12201 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# V_LOW -0.00665f
C12202 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.87e-19
C12203 FALLING_COUNTER.COUNT_SUB_DFF14.Q V_LOW 2.25f
C12204 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# sky130_fd_sc_hd__conb_1_47/HI 5.11e-19
C12205 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__inv_1_30/Y 4.33e-19
C12206 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# -0.00592f
C12207 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 5.25e-21
C12208 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# -4.66e-20
C12209 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__conb_1_17/HI 6.12e-19
C12210 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.97e-19
C12211 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 3.02e-19
C12212 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__conb_1_12/HI 0.0188f
C12213 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.00516f
C12214 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.00346f
C12215 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# -0.0659f
C12216 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__inv_1_39/Y 8.87e-19
C12217 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0488f
C12218 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_64/Y 0.00686f
C12219 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.26e-20
C12220 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__conb_1_16/HI -6.57e-19
C12221 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# -1.44e-20
C12222 sky130_fd_sc_hd__conb_1_10/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 1.2e-19
C12223 sky130_fd_sc_hd__nand3_1_1/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.56e-19
C12224 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__inv_1_41/Y 1.07e-20
C12225 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_5/HI 2.3e-21
C12226 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_1_44/A 0.0209f
C12227 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__conb_1_8/HI 0.00226f
C12228 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# -0.0193f
C12229 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 1.53e-21
C12230 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__conb_1_23/HI 0.0229f
C12231 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_19/HI 3.07e-21
C12232 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_66/A 1.16e-19
C12233 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 0.00189f
C12234 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 1.92e-20
C12235 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# -3.46e-20
C12236 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__conb_1_17/HI 0.103f
C12237 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0233f
C12238 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0156f
C12239 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__conb_1_27/HI 0.0073f
C12240 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__conb_1_34/HI -0.0111f
C12241 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_38/HI 4.32e-19
C12242 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_44/Y 1.24f
C12243 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 6.36e-19
C12244 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__conb_1_20/HI 3.27e-21
C12245 sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 0.254f
C12246 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 7.44e-20
C12247 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__inv_1_40/Y 0.0036f
C12248 FULL_COUNTER.COUNT_SUB_DFF2.Q V_HIGH 0.848f
C12249 sky130_fd_sc_hd__conb_1_25/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.144f
C12250 sky130_fd_sc_hd__inv_1_46/A V_LOW 0.639f
C12251 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_941_21# -0.00122f
C12252 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# -2.3e-19
C12253 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00807f
C12254 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 6.25e-20
C12255 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# -0.00591f
C12256 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# -0.00631f
C12257 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0138f
C12258 sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0335f
C12259 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.0212f
C12260 sky130_fd_sc_hd__conb_1_32/HI V_LOW 0.155f
C12261 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 9.13e-20
C12262 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 7.44e-19
C12263 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00226f
C12264 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_1_29/Y 7.95e-22
C12265 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__inv_1_28/Y 3.76e-21
C12266 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 7.44e-20
C12267 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_34/LO 0.00142f
C12268 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 7.26e-19
C12269 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__conb_1_10/HI 7.32e-19
C12270 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.2e-19
C12271 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00157f
C12272 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.22e-19
C12273 FULL_COUNTER.COUNT_SUB_DFF4.Q V_LOW 0.533f
C12274 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_16_4/Y 7.7e-20
C12275 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_44/Y 1.79f
C12276 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 7.48e-20
C12277 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI -9.25e-19
C12278 V_SENSE FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0036f
C12279 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__inv_1_38/Y 0.0463f
C12280 V_SENSE sky130_fd_sc_hd__inv_16_28/Y 0.0323f
C12281 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_31/HI 2.43e-20
C12282 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__conb_1_16/HI 1.46e-20
C12283 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 3.33e-19
C12284 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# -0.00141f
C12285 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.00558f
C12286 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 1.01e-20
C12287 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0.00523f
C12288 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 9.21e-20
C12289 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# V_LOW -1.39e-35
C12290 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_32/HI 0.0392f
C12291 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00151f
C12292 sky130_fd_sc_hd__conb_1_25/HI FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.47e-19
C12293 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_27/Y 0.0051f
C12294 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 7.91e-20
C12295 sky130_fd_sc_hd__inv_16_51/A CLOCK_GEN.SR_Op.Q 0.0271f
C12296 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 8.96e-19
C12297 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_16_19/Y 2.72e-19
C12298 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__conb_1_12/HI 0.00257f
C12299 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# V_LOW 4.8e-20
C12300 sky130_fd_sc_hd__inv_1_69/Y V_LOW 0.424f
C12301 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__conb_1_4/HI 0.00427f
C12302 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00242f
C12303 sky130_fd_sc_hd__inv_16_41/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0292f
C12304 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_47/Y 0.0956f
C12305 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.0224f
C12306 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.00132f
C12307 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00113f
C12308 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_23/Y 0.0213f
C12309 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -5.54e-21
C12310 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.78e-21
C12311 sky130_fd_sc_hd__inv_1_68/Y V_LOW 0.175f
C12312 FALLING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0727f
C12313 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# V_LOW 1.38e-19
C12314 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__nand2_8_0/a_27_47# 0.022f
C12315 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.52e-19
C12316 sky130_fd_sc_hd__inv_1_24/A V_LOW 0.488f
C12317 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 4.76e-19
C12318 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 1.38e-20
C12319 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 5.32e-20
C12320 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 2.42e-20
C12321 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 8.26e-20
C12322 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00102f
C12323 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# sky130_fd_sc_hd__inv_1_25/Y 7.05e-19
C12324 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__conb_1_38/HI 0.00197f
C12325 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 2.45e-19
C12326 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 6.82e-20
C12327 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_64/Y 0.0813f
C12328 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# 1.19e-19
C12329 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_41/Y 9.8e-20
C12330 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# V_LOW 0.00256f
C12331 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_45/LO 0.0724f
C12332 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# -1.65e-19
C12333 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# -0.00389f
C12334 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# -0.0103f
C12335 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 3.08e-19
C12336 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00203f
C12337 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00178f
C12338 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__inv_1_7/Y 0.00784f
C12339 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0.0011f
C12340 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0662f
C12341 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_49/Y 3.89e-20
C12342 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_67/A 0.00165f
C12343 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 0.0171f
C12344 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# V_LOW 3.56e-20
C12345 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 1.63e-20
C12346 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__conb_1_39/LO 2.12e-19
C12347 sky130_fd_sc_hd__dfbbn_1_28/Q_N RISING_COUNTER.COUNT_SUB_DFF8.Q 0.0069f
C12348 sky130_fd_sc_hd__nand2_8_4/Y sky130_fd_sc_hd__inv_1_66/Y 8.77e-22
C12349 sky130_fd_sc_hd__inv_1_66/Y Reset 0.00856f
C12350 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 4.74e-21
C12351 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0495f
C12352 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 1.13e-20
C12353 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.18e-20
C12354 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__conb_1_51/HI 8.26e-19
C12355 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__conb_1_12/HI 0.00576f
C12356 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__conb_1_24/HI 6.08e-21
C12357 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.109f
C12358 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 2.57e-21
C12359 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 0.00113f
C12360 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 2.69e-19
C12361 sky130_fd_sc_hd__inv_1_51/Y CLOCK_GEN.SR_Op.Q 0.0114f
C12362 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.0113f
C12363 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_56/A 0.00365f
C12364 sky130_fd_sc_hd__nand3_1_1/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 2.47e-20
C12365 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_647_21# -0.00504f
C12366 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# V_LOW 4.8e-20
C12367 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_10/HI -3.44e-19
C12368 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 4.66e-19
C12369 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.00106f
C12370 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 0.00122f
C12371 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 5.05e-19
C12372 FALLING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 2.53e-19
C12373 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__conb_1_29/HI -1.06e-20
C12374 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 6.4e-20
C12375 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.44e-19
C12376 sky130_fd_sc_hd__conb_1_35/HI Reset 0.0389f
C12377 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00636f
C12378 sky130_fd_sc_hd__dfbbn_1_34/Q_N V_LOW -0.0104f
C12379 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_50/Y 0.0519f
C12380 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__conb_1_26/HI 2.06e-20
C12381 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00157f
C12382 sky130_fd_sc_hd__inv_1_39/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00964f
C12383 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_33/Y 0.127f
C12384 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_67/A 0.0498f
C12385 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.42e-19
C12386 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__conb_1_44/HI 0.0108f
C12387 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_1_35/Y 3.08e-20
C12388 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# -8.23e-19
C12389 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# -0.00834f
C12390 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0403f
C12391 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00472f
C12392 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 1.67e-21
C12393 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__nand2_8_4/Y 0.00193f
C12394 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# Reset 0.00718f
C12395 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# -0.00228f
C12396 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# -4.84e-19
C12397 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_24/Y 0.287f
C12398 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_28/Y 9.42e-19
C12399 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__conb_1_4/HI 2.17e-19
C12400 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_24/Y 1.69e-19
C12401 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__conb_1_37/HI 0.00181f
C12402 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00529f
C12403 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# 2.44e-19
C12404 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 4.3e-19
C12405 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 3.04e-19
C12406 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 4.36e-19
C12407 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# -0.00122f
C12408 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# -2.52e-19
C12409 sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__conb_1_30/HI 0.0345f
C12410 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_1_41/Y 5.85e-22
C12411 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_46/HI 0.00207f
C12412 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_17/LO 5.31e-19
C12413 sky130_fd_sc_hd__inv_1_50/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.224f
C12414 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 5.65e-20
C12415 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# 3.67e-21
C12416 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 8e-21
C12417 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 3.28e-20
C12418 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_891_329# 1.97e-20
C12419 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00296f
C12420 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_791_47# 2.82e-19
C12421 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__inv_1_12/Y 2.81e-20
C12422 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.0107f
C12423 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# -6.43e-20
C12424 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# -0.00988f
C12425 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0.0387f
C12426 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# V_LOW 0.0178f
C12427 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# sky130_fd_sc_hd__inv_16_41/Y 6.95e-21
C12428 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# V_LOW 3.56e-20
C12429 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__conb_1_46/HI 2.6e-19
C12430 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__conb_1_18/HI 1.04e-19
C12431 FULL_COUNTER.COUNT_SUB_DFF5.Q V_LOW 0.828f
C12432 sky130_fd_sc_hd__conb_1_47/LO sky130_fd_sc_hd__conb_1_47/HI 0.00538f
C12433 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nor2_1_0/Y 0.00103f
C12434 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# -6.8e-19
C12435 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -0.00453f
C12436 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__inv_1_12/Y 7.31e-19
C12437 sky130_fd_sc_hd__dfbbn_1_31/Q_N RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00254f
C12438 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# RISING_COUNTER.COUNT_SUB_DFF8.Q 9.3e-19
C12439 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# -0.00486f
C12440 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_891_329# -0.00159f
C12441 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 6.43e-20
C12442 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 0.0199f
C12443 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.0148f
C12444 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_53/Y 6.99e-20
C12445 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# V_LOW -0.00121f
C12446 sky130_fd_sc_hd__conb_1_24/LO FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0504f
C12447 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.74e-21
C12448 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF2.Q 2.22e-21
C12449 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_1_7/Y 0.0014f
C12450 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 9.77e-19
C12451 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 2.26e-21
C12452 FULL_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.742f
C12453 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 4.43e-21
C12454 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00313f
C12455 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00595f
C12456 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 0.789f
C12457 sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# sky130_fd_sc_hd__conb_1_12/HI 2.09e-19
C12458 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.319f
C12459 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# sky130_fd_sc_hd__inv_1_37/Y 3.36e-19
C12460 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 2.65e-20
C12461 sky130_fd_sc_hd__inv_1_7/Y V_LOW 0.133f
C12462 sky130_fd_sc_hd__conb_1_18/HI RISING_COUNTER.COUNT_SUB_DFF15.Q 0.115f
C12463 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__conb_1_32/HI 3.77e-19
C12464 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 0.0112f
C12465 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_581_47# -2.6e-20
C12466 sky130_fd_sc_hd__inv_16_19/Y CLOCK_GEN.SR_Op.Q 3.85e-21
C12467 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.00109f
C12468 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_29/Q_N 0.0059f
C12469 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 4.17e-20
C12470 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# sky130_fd_sc_hd__conb_1_29/HI -2.92e-20
C12471 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 7.41e-19
C12472 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 4.18e-19
C12473 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0273f
C12474 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_50/HI 3.1e-20
C12475 sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# sky130_fd_sc_hd__conb_1_26/HI 1.06e-19
C12476 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__inv_1_50/Y 1.72e-20
C12477 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__conb_1_50/HI 2.46e-20
C12478 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 1.04e-19
C12479 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 1.75e-20
C12480 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# -0.00151f
C12481 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# -2.47e-19
C12482 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0012f
C12483 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__conb_1_16/HI 8.83e-21
C12484 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# sky130_fd_sc_hd__conb_1_43/HI 0.00115f
C12485 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0164f
C12486 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__nand2_8_4/Y 1.32e-19
C12487 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# Reset 0.00273f
C12488 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# -9.32e-20
C12489 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_16_41/Y 0.145f
C12490 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# CLOCK_GEN.SR_Op.Q 7.9e-19
C12491 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__conb_1_37/HI 0.00335f
C12492 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.32e-20
C12493 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0216f
C12494 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# -1.76e-19
C12495 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# -0.00115f
C12496 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0359f
C12497 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 7.82e-20
C12498 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/Q_N -4.78e-20
C12499 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__conb_1_29/LO 5.58e-20
C12500 sky130_fd_sc_hd__inv_1_59/Y V_LOW 0.22f
C12501 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.184f
C12502 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0.00107f
C12503 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.108f
C12504 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__inv_1_36/Y 1.31e-20
C12505 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# -9.88e-20
C12506 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -6.23e-21
C12507 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# -0.00367f
C12508 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00113f
C12509 sky130_fd_sc_hd__dfbbn_1_51/Q_N FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00177f
C12510 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__conb_1_4/HI 3.98e-20
C12511 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_0/HI 0.00574f
C12512 sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__conb_1_40/HI 0.00239f
C12513 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_44/A 2.21e-19
C12514 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.00709f
C12515 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# V_LOW -6.55e-19
C12516 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_647_21# -0.00119f
C12517 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__conb_1_46/HI -0.0097f
C12518 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__conb_1_18/HI 9.37e-21
C12519 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_47/Y 4.33e-21
C12520 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 7.19e-19
C12521 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00147f
C12522 sky130_fd_sc_hd__dfbbn_1_40/Q_N V_LOW -2.68e-19
C12523 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# V_LOW 4.8e-20
C12524 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 0.00122f
C12525 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# 3.48e-20
C12526 sky130_fd_sc_hd__nand2_8_9/A FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00182f
C12527 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 7.85e-20
C12528 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_21/LO 3.04e-20
C12529 sky130_fd_sc_hd__nand2_8_8/A CLOCK_GEN.SR_Op.Q 0.0066f
C12530 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_22/Y 1.29e-19
C12531 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# -2.52e-19
C12532 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -4.39e-19
C12533 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 5.65e-20
C12534 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__conb_1_9/HI 8.37e-19
C12535 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# -3.46e-20
C12536 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# V_LOW 2.26e-20
C12537 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00292f
C12538 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 0.00113f
C12539 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_1_44/A 0.00742f
C12540 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.00169f
C12541 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_32/HI 0.0031f
C12542 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_5/HI -0.0148f
C12543 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__conb_1_7/HI 0.00329f
C12544 sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_16_24/Y 0.00203f
C12545 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 9.8e-20
C12546 sky130_fd_sc_hd__dfbbn_1_33/Q_N RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0163f
C12547 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 3e-21
C12548 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_1_44/A 0.0119f
C12549 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00246f
C12550 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_21/Y 0.225f
C12551 sky130_fd_sc_hd__inv_4_0/A FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0025f
C12552 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_1_13/Y 1.2e-20
C12553 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__conb_1_32/HI 0.00262f
C12554 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_20/Y 4.42e-19
C12555 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# V_LOW 4.8e-20
C12556 sky130_fd_sc_hd__inv_1_9/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 3.16e-20
C12557 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 0.00942f
C12558 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# -0.00717f
C12559 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_557_413# -3.67e-20
C12560 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__conb_1_25/HI 0.0037f
C12561 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 5.13e-19
C12562 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__inv_1_13/Y 1.92e-20
C12563 sky130_fd_sc_hd__dfbbn_1_0/Q_N FULL_COUNTER.COUNT_SUB_DFF5.Q 0.021f
C12564 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.78e-19
C12565 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 1.51e-19
C12566 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 7.22e-20
C12567 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__conb_1_35/HI 1.07e-21
C12568 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# 0.00226f
C12569 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 1.89e-20
C12570 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# V_LOW 0.0381f
C12571 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# -7.17e-20
C12572 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# -1.76e-19
C12573 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0268f
C12574 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# V_LOW 0.0122f
C12575 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__inv_1_59/Y 0.0037f
C12576 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 0.0102f
C12577 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/Q_N -9.56e-20
C12578 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_1_64/Y 0.0105f
C12579 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/Q_N 9.65e-21
C12580 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/Q_N -4.78e-20
C12581 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# V_LOW 0.00566f
C12582 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.69e-19
C12583 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.03e-19
C12584 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 7.05e-19
C12585 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_26/Y 2.07e-20
C12586 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__conb_1_37/HI 0.0155f
C12587 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.341f
C12588 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0031f
C12589 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.92e-21
C12590 sky130_fd_sc_hd__inv_16_49/Y sky130_fd_sc_hd__inv_16_50/A 0.932f
C12591 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 2.25e-21
C12592 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 9.42e-20
C12593 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0052f
C12594 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# -2.07e-19
C12595 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0603f
C12596 sky130_fd_sc_hd__nand2_1_1/a_113_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.9e-19
C12597 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# V_LOW 0.00829f
C12598 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__conb_1_33/HI -3.29e-19
C12599 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__conb_1_2/HI 3.85e-21
C12600 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__conb_1_12/HI 6.29e-19
C12601 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 0.00157f
C12602 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.012f
C12603 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 6.1e-21
C12604 RISING_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.277f
C12605 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.014f
C12606 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 0.0124f
C12607 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 5.69e-20
C12608 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# -0.00753f
C12609 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.00244f
C12610 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 0.0174f
C12611 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__inv_1_69/Y 0.00243f
C12612 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 6.47e-19
C12613 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0294f
C12614 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_1_60/Y 0.16f
C12615 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_581_47# -2.6e-20
C12616 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_67/A 6.28e-20
C12617 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 9.07e-19
C12618 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.48e-19
C12619 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# V_LOW 0.00942f
C12620 sky130_fd_sc_hd__inv_1_8/Y V_LOW 0.295f
C12621 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/Q_N 8.96e-21
C12622 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0136f
C12623 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# sky130_fd_sc_hd__inv_1_22/Y 1.69e-19
C12624 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 3.54e-21
C12625 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# sky130_fd_sc_hd__conb_1_28/HI 8.26e-19
C12626 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__conb_1_5/HI 2.87e-20
C12627 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# -1.76e-19
C12628 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# -7.17e-20
C12629 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_16_41/Y 4.02e-19
C12630 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.78e-20
C12631 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 0.0327f
C12632 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__conb_1_32/HI 0.00103f
C12633 sky130_fd_sc_hd__nand2_8_9/a_27_47# V_LOW -0.0117f
C12634 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.04e-20
C12635 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# sky130_fd_sc_hd__conb_1_5/HI 4.85e-19
C12636 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.0124f
C12637 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.00799f
C12638 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 6.02e-19
C12639 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0395f
C12640 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__inv_1_2/Y 2.87e-20
C12641 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_20/HI 8.37e-20
C12642 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_49/Y 5.19e-20
C12643 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_1_44/A 1.32e-21
C12644 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.175f
C12645 sky130_fd_sc_hd__inv_1_38/Y sky130_fd_sc_hd__conb_1_30/HI 0.165f
C12646 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 4.22e-21
C12647 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00211f
C12648 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# -0.00522f
C12649 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# 0.00111f
C12650 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__conb_1_17/HI 0.0175f
C12651 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# 2.06e-20
C12652 FALLING_COUNTER.COUNT_SUB_DFF0.Q V_LOW 1.53f
C12653 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__conb_1_30/HI 0.0132f
C12654 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00206f
C12655 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# sky130_fd_sc_hd__conb_1_25/HI 2.78e-21
C12656 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.00157f
C12657 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__conb_1_8/LO 5.88e-22
C12658 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_1_39/Y 3.06e-19
C12659 sky130_fd_sc_hd__inv_16_16/Y V_LOW 0.161f
C12660 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_381_47# 0.014f
C12661 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__conb_1_0/HI 0.0203f
C12662 sky130_fd_sc_hd__inv_1_58/Y V_LOW 0.025f
C12663 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 0.0348f
C12664 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# V_LOW 2.94e-20
C12665 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__conb_1_45/HI 0.0431f
C12666 sky130_fd_sc_hd__conb_1_50/HI RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0242f
C12667 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00135f
C12668 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# V_LOW 4.7e-20
C12669 V_SENSE sky130_fd_sc_hd__inv_16_20/A 0.00314f
C12670 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0.00316f
C12671 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__conb_1_37/HI 4.3e-21
C12672 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 9.68e-20
C12673 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_23/HI 2.08e-21
C12674 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_64/Y 0.0838f
C12675 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__conb_1_7/LO 0.134f
C12676 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.00121f
C12677 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# V_LOW 0.00351f
C12678 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__conb_1_11/HI 3.33e-21
C12679 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 6.45e-21
C12680 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 5.18e-20
C12681 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 4.97e-19
C12682 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_16_4/Y 1.32e-19
C12683 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00654f
C12684 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0192f
C12685 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_10/Y 0.333f
C12686 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.00212f
C12687 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_6/HI 0.00398f
C12688 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# V_LOW 3.56e-20
C12689 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# -3.86e-20
C12690 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# -1.61e-20
C12691 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# 8.48e-19
C12692 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__conb_1_12/HI 6.52e-20
C12693 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00715f
C12694 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__conb_1_37/HI 2.86e-19
C12695 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_7/HI 6.64e-21
C12696 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# 7.12e-19
C12697 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_581_47# 4.18e-19
C12698 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# -0.00141f
C12699 sky130_fd_sc_hd__inv_2_0/A FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0186f
C12700 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__conb_1_31/HI 0.00101f
C12701 sky130_fd_sc_hd__nand2_8_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.06e-19
C12702 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_11/LO 9.95e-20
C12703 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0348f
C12704 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_1_41/Y 6.11e-20
C12705 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.53e-19
C12706 sky130_fd_sc_hd__dfbbn_1_50/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 5.62e-20
C12707 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_1_5/Y 0.0416f
C12708 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.11e-19
C12709 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.92e-22
C12710 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# V_LOW 1.79e-20
C12711 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.012f
C12712 sky130_fd_sc_hd__nand3_1_2/a_109_47# CLOCK_GEN.SR_Op.Q 6.25e-19
C12713 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_557_413# -3.67e-20
C12714 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# -0.00623f
C12715 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__conb_1_21/LO 3.08e-19
C12716 sky130_fd_sc_hd__inv_16_16/Y sky130_fd_sc_hd__inv_16_9/Y 2.13e-19
C12717 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0234f
C12718 sky130_fd_sc_hd__dfbbn_1_19/a_1159_47# sky130_fd_sc_hd__inv_1_25/Y 7.5e-20
C12719 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0161f
C12720 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_791_47# 0.0365f
C12721 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.43e-19
C12722 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF12.Q 1.42e-21
C12723 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_61/Y 3.97e-21
C12724 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__conb_1_2/HI 9.04e-20
C12725 RISING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.81f
C12726 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 2.97e-19
C12727 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__conb_1_47/LO 8.84e-20
C12728 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.0281f
C12729 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 6.34e-19
C12730 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# V_LOW -0.0816f
C12731 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 5.07e-21
C12732 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# Reset 7.19e-19
C12733 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__inv_1_58/Y 0.0025f
C12734 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__inv_1_0/Y 0.132f
C12735 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_25/LO 0.00696f
C12736 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__conb_1_23/HI 9.42e-19
C12737 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_16/a_557_413# 9.02e-19
C12738 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_53/A 4.75e-19
C12739 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF2.Q 3.8e-19
C12740 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_1/Y 0.066f
C12741 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_581_47# -7.91e-19
C12742 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00777f
C12743 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.09e-19
C12744 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 4.24e-19
C12745 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# -3.79e-20
C12746 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# -0.00336f
C12747 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_1_60/Y 0.0409f
C12748 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__conb_1_8/LO 5.59e-20
C12749 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# sky130_fd_sc_hd__inv_1_39/Y 7.69e-22
C12750 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__inv_1_14/Y 0.00188f
C12751 sky130_fd_sc_hd__inv_1_3/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0221f
C12752 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# sky130_fd_sc_hd__conb_1_0/HI 4.96e-20
C12753 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_41/HI 0.00134f
C12754 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# sky130_fd_sc_hd__conb_1_45/HI 4.99e-19
C12755 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0.0225f
C12756 sky130_fd_sc_hd__dfbbn_1_14/Q_N V_LOW -0.00141f
C12757 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_1_19/A 0.0434f
C12758 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 0.00665f
C12759 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.34e-19
C12760 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/Q_N 0.0016f
C12761 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.57e-21
C12762 sky130_fd_sc_hd__inv_1_47/Y CLOCK_GEN.SR_Op.Q 0.675f
C12763 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00187f
C12764 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_6/LO 8.84e-20
C12765 sky130_fd_sc_hd__inv_16_9/A sky130_fd_sc_hd__inv_16_8/A 0.00666f
C12766 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0169f
C12767 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 1.47e-20
C12768 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0114f
C12769 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0.00264f
C12770 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0199f
C12771 sky130_fd_sc_hd__dfbbn_1_47/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.73e-19
C12772 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_29/HI 2.59e-22
C12773 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__conb_1_50/HI 8.72e-19
C12774 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_16_42/Y 2.33e-19
C12775 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.00221f
C12776 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__conb_1_6/HI 3.48e-20
C12777 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/a_941_21# 1.89e-19
C12778 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 8.72e-20
C12779 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 4.27e-19
C12780 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00209f
C12781 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# -2.57e-20
C12782 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__conb_1_12/HI 0.0157f
C12783 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__inv_1_28/Y 6.93e-20
C12784 sky130_fd_sc_hd__dfbbn_1_0/Q_N FALLING_COUNTER.COUNT_SUB_DFF0.Q 4.52e-22
C12785 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_53/Y 4.82e-22
C12786 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# sky130_fd_sc_hd__inv_2_0/A 0.00224f
C12787 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__conb_1_41/HI 7.68e-19
C12788 sky130_fd_sc_hd__inv_1_47/A FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0302f
C12789 sky130_fd_sc_hd__inv_16_22/A sky130_fd_sc_hd__inv_16_8/A 8.42e-20
C12790 sky130_fd_sc_hd__inv_16_29/Y sky130_fd_sc_hd__inv_16_8/Y 0.0152f
C12791 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_1_21/Y 2.68e-19
C12792 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__conb_1_45/HI 1.36e-20
C12793 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_18/A 0.0208f
C12794 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# -3.86e-20
C12795 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# -0.004f
C12796 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0202f
C12797 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_647_21# -0.00889f
C12798 sky130_fd_sc_hd__dfbbn_1_7/Q_N FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00501f
C12799 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00741f
C12800 RISING_COUNTER.COUNT_SUB_DFF0.Q V_LOW 0.856f
C12801 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0482f
C12802 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_51/HI 0.00681f
C12803 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_1_35/Y 3.77e-20
C12804 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 1.12e-20
C12805 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 3.86e-20
C12806 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 2.22e-20
C12807 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_55/Y 0.184f
C12808 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 8e-21
C12809 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 3.67e-21
C12810 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 2.64e-19
C12811 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_24/HI 4.69e-20
C12812 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# V_LOW 2.26e-20
C12813 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__nand2_8_9/A 1.67e-19
C12814 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 3.26e-20
C12815 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 3.71e-19
C12816 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# V_LOW -2.68e-19
C12817 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 4.1e-19
C12818 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 4.56e-20
C12819 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.58e-21
C12820 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# CLOCK_GEN.SR_Op.Q 3.76e-21
C12821 sky130_fd_sc_hd__inv_16_4/Y Reset 1.68e-19
C12822 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_24/HI 0.0237f
C12823 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# V_LOW 3.56e-20
C12824 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_4_0/A 3.46e-20
C12825 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__conb_1_6/HI 3.44e-19
C12826 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.5e-20
C12827 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00225f
C12828 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00224f
C12829 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00114f
C12830 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 9.52e-20
C12831 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_9/HI 1.59e-19
C12832 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 7.89e-21
C12833 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# -3.79e-20
C12834 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# -4.66e-20
C12835 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# V_LOW 4.8e-20
C12836 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# V_LOW 0.0097f
C12837 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__inv_1_39/Y 0.00421f
C12838 sky130_fd_sc_hd__nand2_8_9/A FULL_COUNTER.COUNT_SUB_DFF0.Q 4.78e-19
C12839 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00194f
C12840 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_67/Y 2.07e-20
C12841 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__inv_1_8/Y 0.00591f
C12842 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 0.00314f
C12843 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.0379f
C12844 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__conb_1_41/HI -0.00686f
C12845 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 0.00525f
C12846 V_SENSE sky130_fd_sc_hd__inv_16_7/A 6.26e-19
C12847 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_47/Y 1.27e-20
C12848 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__inv_1_61/Y 5.54e-19
C12849 sky130_fd_sc_hd__inv_1_41/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0134f
C12850 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# sky130_fd_sc_hd__conb_1_4/HI 4.94e-19
C12851 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0187f
C12852 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 8.44e-20
C12853 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 2.4e-19
C12854 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# sky130_fd_sc_hd__conb_1_19/HI 4.7e-20
C12855 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__conb_1_29/HI 8.67e-20
C12856 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.0245f
C12857 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__conb_1_41/HI 8.84e-20
C12858 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__conb_1_26/HI 2.52e-19
C12859 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_891_329# -2.2e-20
C12860 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# -4.1e-19
C12861 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__conb_1_6/HI 8.96e-21
C12862 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_16/LO 1.14e-19
C12863 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_32/Y 0.0177f
C12864 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 6.42e-21
C12865 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__conb_1_51/HI 5.23e-19
C12866 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/Q_N 4.28e-21
C12867 sky130_fd_sc_hd__inv_1_43/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 8.03e-21
C12868 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# sky130_fd_sc_hd__conb_1_47/HI 0.00286f
C12869 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00256f
C12870 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 1.48e-20
C12871 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 4.49e-20
C12872 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__conb_1_51/HI 0.00282f
C12873 sky130_fd_sc_hd__inv_1_9/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 7.54e-21
C12874 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__conb_1_15/LO 2.41e-20
C12875 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_647_21# -0.00548f
C12876 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.00669f
C12877 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__inv_1_31/Y 4.56e-21
C12878 sky130_fd_sc_hd__nand2_1_2/a_113_47# V_LOW -1.78e-19
C12879 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# Reset 2.24e-21
C12880 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# sky130_fd_sc_hd__inv_1_44/A 7.83e-19
C12881 sky130_fd_sc_hd__conb_1_16/HI FULL_COUNTER.COUNT_SUB_DFF16.Q 1.62e-19
C12882 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00586f
C12883 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__conb_1_25/LO 1.31e-20
C12884 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# -8.41e-19
C12885 sky130_fd_sc_hd__conb_1_35/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00249f
C12886 sky130_fd_sc_hd__inv_1_57/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00457f
C12887 FALLING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.974f
C12888 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 0.0243f
C12889 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__conb_1_15/HI 0.00771f
C12890 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 4.16e-19
C12891 sky130_fd_sc_hd__conb_1_43/HI V_LOW 0.104f
C12892 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_581_47# -2.6e-20
C12893 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0425f
C12894 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__conb_1_25/HI 1.36e-20
C12895 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0165f
C12896 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 1.44e-20
C12897 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# sky130_fd_sc_hd__inv_1_55/Y 2.59e-19
C12898 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__inv_1_33/Y 2.02e-19
C12899 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__conb_1_15/HI -8.28e-19
C12900 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__conb_1_11/HI 1.24e-19
C12901 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__conb_1_8/HI 3.87e-19
C12902 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# -0.0122f
C12903 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -4.52e-19
C12904 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 2.2e-20
C12905 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# V_LOW 0.0124f
C12906 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 6.6e-19
C12907 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# V_LOW -0.00266f
C12908 sky130_fd_sc_hd__nand2_8_4/a_27_47# CLOCK_GEN.SR_Op.Q 0.0384f
C12909 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# -4.66e-20
C12910 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# -6.94e-36
C12911 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# V_LOW -0.324f
C12912 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 2.13f
C12913 sky130_fd_sc_hd__inv_8_0/A FULL_COUNTER.COUNT_SUB_DFF0.Q 2.15e-20
C12914 sky130_fd_sc_hd__conb_1_3/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 5.15e-21
C12915 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_56/Y 2.98e-19
C12916 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.22e-20
C12917 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# V_LOW -0.00266f
C12918 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.5e-19
C12919 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# V_LOW 2.66e-19
C12920 sky130_fd_sc_hd__dfbbn_1_47/a_581_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 7.56e-20
C12921 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q -5.81e-37
C12922 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__conb_1_7/HI 0.00571f
C12923 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# V_LOW 0.00877f
C12924 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_42/LO 9.32e-20
C12925 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# sky130_fd_sc_hd__inv_16_41/Y 8.68e-19
C12926 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 0.0112f
C12927 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# V_LOW -0.00268f
C12928 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# V_LOW -1.01e-19
C12929 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_24/Y 5.9e-22
C12930 sky130_fd_sc_hd__dfbbn_1_0/Q_N RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0169f
C12931 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.0416f
C12932 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_13/LO 9.74e-21
C12933 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__nand2_8_9/A 9.18e-19
C12934 V_SENSE sky130_fd_sc_hd__inv_1_50/Y 1.59e-19
C12935 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_7/HI 3.8e-20
C12936 sky130_fd_sc_hd__inv_16_41/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.288f
C12937 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_42/Y 7.12e-20
C12938 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0339f
C12939 sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 1.52f
C12940 sky130_fd_sc_hd__conb_1_27/LO FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0132f
C12941 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 1.68e-19
C12942 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 0.317f
C12943 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__conb_1_29/HI 1.69e-19
C12944 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_5/HI 8.15e-19
C12945 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# V_LOW -0.313f
C12946 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1_19/Y 0.00207f
C12947 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# V_LOW 1.38e-19
C12948 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__conb_1_26/HI 2.43e-19
C12949 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# -1.42e-32
C12950 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# -0.00385f
C12951 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.6e-20
C12952 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 8.99e-20
C12953 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 1.07e-20
C12954 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__conb_1_51/HI 0.00215f
C12955 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.37e-20
C12956 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__conb_1_44/HI 0.0179f
C12957 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.097f
C12958 FULL_COUNTER.COUNT_SUB_DFF1.Q V_LOW 2.14f
C12959 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_581_47# -2.6e-20
C12960 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__inv_1_41/Y 5.89e-21
C12961 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_3/a_941_21# -5.45e-20
C12962 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.00207f
C12963 sky130_fd_sc_hd__inv_16_4/Y sky130_fd_sc_hd__inv_1_44/A 0.0077f
C12964 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 0.0202f
C12965 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# V_LOW -0.00121f
C12966 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_8_0/A 6.98e-20
C12967 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__conb_1_49/LO 4.83e-20
C12968 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# sky130_fd_sc_hd__conb_1_6/HI 3.15e-19
C12969 sky130_fd_sc_hd__conb_1_50/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.44e-19
C12970 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__conb_1_15/HI 4.06e-19
C12971 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 4.42e-20
C12972 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 4.42e-20
C12973 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 7.69e-20
C12974 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.64e-19
C12975 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 6.97e-22
C12976 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__inv_16_40/Y 0.431f
C12977 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__inv_1_33/Y 5.95e-21
C12978 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 2.59e-19
C12979 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__conb_1_15/HI -2.07e-19
C12980 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 8.88e-20
C12981 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 3.38e-19
C12982 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__conb_1_33/HI 2.67e-20
C12983 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# 0.00138f
C12984 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__conb_1_8/HI -0.01f
C12985 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_6/HI 0.00185f
C12986 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 1.54e-22
C12987 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.26e-20
C12988 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# -2.37e-19
C12989 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -0.00447f
C12990 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# -2.57e-20
C12991 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.38e-20
C12992 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_20/HI 4.67e-19
C12993 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_17/HI 7.81e-19
C12994 sky130_fd_sc_hd__inv_2_0/A FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0981f
C12995 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_647_21# -0.00631f
C12996 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_473_413# -0.0147f
C12997 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 1.47e-21
C12998 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.62e-19
C12999 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# sky130_fd_sc_hd__conb_1_7/HI -8.7e-21
C13000 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00757f
C13001 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# V_LOW 2.94e-20
C13002 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_23/LO 0.0181f
C13003 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# 0.0024f
C13004 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 0.0571f
C13005 sky130_fd_sc_hd__inv_1_43/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00369f
C13006 V_HIGH FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.71f
C13007 FALLING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 9.15e-21
C13008 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__conb_1_40/HI 0.00926f
C13009 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0152f
C13010 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.041f
C13011 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 5.69e-21
C13012 sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0236f
C13013 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__conb_1_24/HI 0.0151f
C13014 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_53/A 0.243f
C13015 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_48/Y 0.00415f
C13016 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00706f
C13017 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__inv_1_13/Y 0.0163f
C13018 sky130_fd_sc_hd__inv_16_44/A sky130_fd_sc_hd__inv_16_55/A 0.0322f
C13019 sky130_fd_sc_hd__inv_16_29/Y sky130_fd_sc_hd__inv_16_29/A 0.0693f
C13020 sky130_fd_sc_hd__inv_1_36/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0768f
C13021 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 2.51f
C13022 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1_15/HI 0.0357f
C13023 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_7/HI 1.17e-19
C13024 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -0.0116f
C13025 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# -2.37e-19
C13026 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0327f
C13027 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 7.25e-19
C13028 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__conb_1_8/HI 0.0116f
C13029 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__conb_1_29/HI 0.00203f
C13030 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 0.00451f
C13031 sky130_fd_sc_hd__fill_8_932/VPB V_LOW 0.797f
C13032 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__conb_1_26/HI 4.38e-20
C13033 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_29/Y 0.015f
C13034 sky130_fd_sc_hd__conb_1_25/HI FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00481f
C13035 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_16_24/Y 7.38e-22
C13036 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_16_40/Y 1.63e-20
C13037 sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__conb_1_32/HI 0.00162f
C13038 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_22/Y 4.83e-19
C13039 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 2.17e-19
C13040 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.021f
C13041 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.58e-19
C13042 sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.203f
C13043 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 6.25e-21
C13044 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_24/HI 7.59e-20
C13045 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__conb_1_44/HI 0.00613f
C13046 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00148f
C13047 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_47/A 3.3e-19
C13048 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# V_LOW -9.15e-19
C13049 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__conb_1_48/HI 0.0106f
C13050 sky130_fd_sc_hd__inv_16_19/Y sky130_fd_sc_hd__inv_1_23/Y 0.00183f
C13051 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.86e-19
C13052 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.06e-19
C13053 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.46e-20
C13054 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00268f
C13055 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0245f
C13056 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.0183f
C13057 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_66/A 0.00493f
C13058 sky130_fd_sc_hd__inv_16_45/A sky130_fd_sc_hd__inv_16_55/A 0.266f
C13059 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__inv_16_42/Y 0.0353f
C13060 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 5.57e-21
C13061 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 0.0397f
C13062 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__inv_1_31/Y 1.36e-20
C13063 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 0.026f
C13064 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 1.45e-19
C13065 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 1.45e-19
C13066 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_2_0/A 0.00202f
C13067 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.028f
C13068 sky130_fd_sc_hd__dfbbn_1_1/Q_N FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0286f
C13069 sky130_fd_sc_hd__conb_1_3/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00665f
C13070 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_193_47# -0.11f
C13071 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.00249f
C13072 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__inv_1_0/Y 0.0388f
C13073 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 0.014f
C13074 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# V_LOW -0.0146f
C13075 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.78e-19
C13076 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__conb_1_10/HI 4.38e-20
C13077 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# -9.35e-20
C13078 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# -3.86e-20
C13079 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_23/Y 0.0164f
C13080 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__conb_1_24/HI 5.37e-19
C13081 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# -1.66e-19
C13082 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_791_47# -2.22e-34
C13083 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 3.21e-20
C13084 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 3.21e-19
C13085 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_10/Y 0.266f
C13086 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_31/Y 8.59e-21
C13087 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__conb_1_35/HI 0.00245f
C13088 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_6/Q_N 3.34e-19
C13089 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.25e-20
C13090 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__conb_1_40/HI 0.00613f
C13091 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 2.72e-20
C13092 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__conb_1_17/HI 9.91e-20
C13093 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.00263f
C13094 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_46/HI 7.38e-20
C13095 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# V_LOW 0.00534f
C13096 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 0.00384f
C13097 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 0.00136f
C13098 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 4.17e-20
C13099 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 8.67e-19
C13100 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# -0.00263f
C13101 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# -5.54e-21
C13102 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 2.36e-21
C13103 RISING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0333f
C13104 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# 0.0037f
C13105 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 2.74e-21
C13106 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_20/HI 4.91e-19
C13107 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.00109f
C13108 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 2.12e-19
C13109 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0016f
C13110 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00621f
C13111 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 9.48e-20
C13112 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 9.48e-20
C13113 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_1_1/Y 0.00331f
C13114 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_2_0/A 1.17e-20
C13115 sky130_fd_sc_hd__dfbbn_1_13/Q_N V_LOW -0.0104f
C13116 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF15.Q 0.014f
C13117 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_8/Y 0.0179f
C13118 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 0.00987f
C13119 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 0.0101f
C13120 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_26/Y 0.0267f
C13121 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.0608f
C13122 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00187f
C13123 sky130_fd_sc_hd__conb_1_16/HI FULL_COUNTER.COUNT_SUB_DFF17.Q 6.17e-20
C13124 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 6.37e-19
C13125 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 4.37e-19
C13126 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.00167f
C13127 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.13e-20
C13128 sky130_fd_sc_hd__inv_16_55/Y sky130_fd_sc_hd__inv_16_50/A 0.00277f
C13129 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# V_LOW -0.102f
C13130 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__conb_1_19/LO 1.47e-20
C13131 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0366f
C13132 FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0111f
C13133 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__conb_1_9/HI 1.62e-20
C13134 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# -1.66e-19
C13135 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# -7.17e-20
C13136 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00493f
C13137 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 1.67e-19
C13138 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# -0.00913f
C13139 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_891_329# -2.2e-20
C13140 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 1.18e-19
C13141 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 9.29e-19
C13142 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0605f
C13143 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 4.13e-20
C13144 sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__inv_1_66/Y 0.00101f
C13145 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.53e-19
C13146 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0064f
C13147 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 7.69e-20
C13148 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__conb_1_14/HI 0.0142f
C13149 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__conb_1_10/HI 0.00771f
C13150 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__conb_1_44/HI 0.00107f
C13151 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__conb_1_48/HI -8.1e-19
C13152 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0482f
C13153 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__conb_1_39/HI 4.86e-20
C13154 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 1.07e-20
C13155 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 1.69e-19
C13156 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__conb_1_35/LO 0.0136f
C13157 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__inv_1_50/Y 4.4e-19
C13158 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__inv_1_14/Y 3.93e-20
C13159 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# -6.57e-19
C13160 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00482f
C13161 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__nand2_8_9/A 0.00243f
C13162 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_0/HI 0.0279f
C13163 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_46/A 0.421f
C13164 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0277f
C13165 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# 2.78e-22
C13166 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00139f
C13167 sky130_fd_sc_hd__inv_1_41/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0221f
C13168 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.15e-20
C13169 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# V_LOW 0.00154f
C13170 sky130_fd_sc_hd__dfbbn_1_46/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 0.00179f
C13171 RISING_COUNTER.COUNT_SUB_DFF0.Q V_HIGH 1.71f
C13172 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# -2.57e-20
C13173 sky130_fd_sc_hd__conb_1_34/LO RISING_COUNTER.COUNT_SUB_DFF8.Q 2.27e-19
C13174 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_0/Y 0.114f
C13175 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 3.19e-19
C13176 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_1_59/Y 0.405f
C13177 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__conb_1_35/HI 0.00213f
C13178 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 4.44e-20
C13179 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 4.33e-22
C13180 sky130_fd_sc_hd__dfbbn_1_38/a_581_47# sky130_fd_sc_hd__conb_1_40/HI 3.73e-19
C13181 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 9.03e-21
C13182 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__conb_1_17/HI 1.96e-19
C13183 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__inv_16_41/Y 0.464f
C13184 sky130_fd_sc_hd__inv_16_28/Y sky130_fd_sc_hd__inv_16_8/A 0.0534f
C13185 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0334f
C13186 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 0.0204f
C13187 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00105f
C13188 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# V_LOW 2.26e-20
C13189 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__inv_16_40/Y 6.2e-21
C13190 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# -0.0592f
C13191 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# -5.78e-20
C13192 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# -0.00631f
C13193 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_1_49/Y 0.00882f
C13194 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0.0262f
C13195 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# 3.78e-19
C13196 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__conb_1_42/LO 9.82e-19
C13197 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# -9.32e-20
C13198 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 1.57e-19
C13199 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# 0.00459f
C13200 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0.00942f
C13201 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# 3.15e-19
C13202 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_24/A 7.96e-19
C13203 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 4.94e-19
C13204 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__conb_1_51/HI 5.29e-19
C13205 sky130_fd_sc_hd__inv_1_57/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 5.37e-20
C13206 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__inv_16_40/Y 0.00187f
C13207 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 7.89f
C13208 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 7.23e-19
C13209 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# 2.65e-20
C13210 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 5.54e-19
C13211 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 1.14e-19
C13212 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00616f
C13213 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_16_41/Y 0.178f
C13214 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.92e-19
C13215 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__inv_1_2/Y 0.00853f
C13216 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# V_LOW 0.0021f
C13217 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__inv_1_30/Y 0.0147f
C13218 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_24/HI 0.0139f
C13219 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_557_413# -3.67e-20
C13220 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# -0.0145f
C13221 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0327f
C13222 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# V_LOW -2.68e-19
C13223 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0429f
C13224 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# sky130_fd_sc_hd__conb_1_9/HI 6.08e-21
C13225 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00383f
C13226 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__conb_1_3/HI -0.00114f
C13227 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# -0.00592f
C13228 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# -1.42e-32
C13229 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__nand3_1_2/Y 1.63e-19
C13230 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.78e-22
C13231 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 6.18e-20
C13232 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF6.Q 2.14e-20
C13233 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# V_LOW 0.0146f
C13234 RISING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00418f
C13235 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 3.11e-22
C13236 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 1.58e-20
C13237 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_1_11/Y 0.00222f
C13238 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__inv_16_42/Y 0.0198f
C13239 sky130_fd_sc_hd__inv_16_44/Y sky130_fd_sc_hd__inv_16_50/A 0.168f
C13240 sky130_fd_sc_hd__dfbbn_1_22/Q_N FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.0285f
C13241 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__conb_1_10/HI 4.06e-19
C13242 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__conb_1_9/HI 7.99e-19
C13243 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__conb_1_48/HI -1.64e-19
C13244 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_9/A 0.00443f
C13245 sky130_fd_sc_hd__inv_1_11/Y V_LOW 0.232f
C13246 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_24/A 0.173f
C13247 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# sky130_fd_sc_hd__conb_1_39/HI 0.00196f
C13248 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.0199f
C13249 sky130_fd_sc_hd__inv_16_40/Y sky130_fd_sc_hd__conb_1_2/HI 0.234f
C13250 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__inv_1_10/Y 0.00128f
C13251 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 9.37e-21
C13252 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0339f
C13253 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_8/LO 3.39e-20
C13254 sky130_fd_sc_hd__inv_1_35/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.122f
C13255 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# Reset 0.00357f
C13256 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_23/HI 0.00252f
C13257 sky130_fd_sc_hd__nand2_1_4/a_113_47# V_LOW -1.78e-19
C13258 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_381_47# 2.26e-21
C13259 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 4.91e-21
C13260 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 5.08e-20
C13261 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 2.42e-20
C13262 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00127f
C13263 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 0.144f
C13264 sky130_fd_sc_hd__conb_1_14/HI V_LOW 0.515f
C13265 sky130_fd_sc_hd__inv_1_3/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 8.78e-20
C13266 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__conb_1_2/HI 3.14e-19
C13267 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00215f
C13268 Reset sky130_fd_sc_hd__conb_1_38/HI 6.45e-21
C13269 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.01e-19
C13270 sky130_fd_sc_hd__conb_1_50/LO RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0161f
C13271 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__inv_1_59/Y 5.77e-20
C13272 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__inv_1_27/Y 8.5e-19
C13273 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__conb_1_29/HI 1.41e-19
C13274 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 4.03e-20
C13275 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_60/Y 9.57e-21
C13276 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF13.Q 1.11e-19
C13277 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.42e-21
C13278 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 0.00114f
C13279 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.05e-20
C13280 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# 0.00226f
C13281 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__inv_1_32/Y 6.38e-20
C13282 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 8.26e-22
C13283 sky130_fd_sc_hd__conb_1_45/HI FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00267f
C13284 sky130_fd_sc_hd__dfbbn_1_9/Q_N V_LOW -0.00141f
C13285 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.96e-19
C13286 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 1.26e-19
C13287 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 1.2e-20
C13288 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# sky130_fd_sc_hd__inv_1_49/Y 2.05e-21
C13289 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0119f
C13290 sky130_fd_sc_hd__nand2_8_5/a_27_47# CLOCK_GEN.SR_Op.Q 7.8e-20
C13291 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/Q_N -4.33e-20
C13292 FULL_COUNTER.COUNT_SUB_DFF0.Q V_LOW 0.708f
C13293 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_1_40/Y 0.00316f
C13294 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_24/Q_N 0.00188f
C13295 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 2.06e-20
C13296 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.94e-19
C13297 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# -0.00263f
C13298 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_891_329# -3.3e-20
C13299 sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__inv_1_38/Y 6.32e-19
C13300 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# sky130_fd_sc_hd__inv_1_3/Y 7.97e-21
C13301 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_40/a_647_21# 7.69e-19
C13302 sky130_fd_sc_hd__conb_1_3/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.22e-21
C13303 sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0738f
C13304 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# 4.17e-19
C13305 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# 2.2e-19
C13306 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.02e-20
C13307 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 2.19e-19
C13308 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.6e-19
C13309 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 2.93e-19
C13310 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0148f
C13311 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 5.08e-20
C13312 sky130_fd_sc_hd__inv_1_32/Y RISING_COUNTER.COUNT_SUB_DFF15.Q 6.94e-20
C13313 FALLING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 2f
C13314 sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__inv_1_59/Y 2.13e-21
C13315 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 2.07e-19
C13316 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# V_LOW 4.61e-20
C13317 sky130_fd_sc_hd__inv_16_2/Y transmission_gate_9/GN 0.0697f
C13318 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# -0.0822f
C13319 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0125f
C13320 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# V_LOW 0.0353f
C13321 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# V_LOW 1.38e-19
C13322 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_16_41/Y 0.321f
C13323 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# -2.53e-20
C13324 sky130_fd_sc_hd__dfbbn_1_48/Q_N FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0063f
C13325 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1_29/LO 1.16e-20
C13326 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0111f
C13327 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 5.21e-21
C13328 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_56/Y 0.096f
C13329 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__conb_1_3/HI -2.07e-19
C13330 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__inv_1_60/Y 5.6e-19
C13331 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.0932f
C13332 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_557_413# -3.67e-20
C13333 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# -0.00279f
C13334 FALLING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 0.768f
C13335 sky130_fd_sc_hd__conb_1_39/HI Reset 0.02f
C13336 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__nand2_8_4/Y 1.26e-19
C13337 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_52/A 2.79e-20
C13338 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# sky130_fd_sc_hd__inv_16_40/Y 0.00297f
C13339 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 4.75e-21
C13340 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# sky130_fd_sc_hd__inv_16_42/Y 0.00118f
C13341 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0302f
C13342 sky130_fd_sc_hd__nor2_1_0/Y CLOCK_GEN.SR_Op.Q 0.121f
C13343 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_891_329# 2.87e-19
C13344 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__inv_1_21/Y 3e-19
C13345 FALLING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 0.64f
C13346 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__conb_1_9/HI 7.22e-19
C13347 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.119f
C13348 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_1_29/Y 0.00101f
C13349 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 0.00117f
C13350 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 8.4e-20
C13351 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 1.48e-20
C13352 V_HIGH FULL_COUNTER.COUNT_SUB_DFF1.Q 1.33f
C13353 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_16_41/Y 0.594f
C13354 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.1e-21
C13355 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.112f
C13356 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 3.45e-19
C13357 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__inv_1_9/Y 1.67e-20
C13358 sky130_fd_sc_hd__inv_16_6/A RISING_COUNTER.COUNT_SUB_DFF4.Q 8.25e-20
C13359 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# sky130_fd_sc_hd__inv_1_27/Y 9.58e-19
C13360 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# Reset 2.28e-19
C13361 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# sky130_fd_sc_hd__conb_1_23/HI 0.00147f
C13362 sky130_fd_sc_hd__inv_1_18/Y V_LOW 0.0315f
C13363 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 2.94e-20
C13364 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# 3.91e-19
C13365 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_1/a_381_47# 8.6e-19
C13366 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.96e-20
C13367 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__inv_16_41/Y 0.0264f
C13368 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 0.0135f
C13369 sky130_fd_sc_hd__inv_1_56/A sky130_fd_sc_hd__inv_1_66/A 0.0786f
C13370 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# sky130_fd_sc_hd__conb_1_2/HI -2.65e-20
C13371 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_0/HI 0.00192f
C13372 sky130_fd_sc_hd__inv_16_7/Y sky130_fd_sc_hd__inv_16_29/A 0.224f
C13373 sky130_fd_sc_hd__dfbbn_1_46/Q_N FALLING_COUNTER.COUNT_SUB_DFF3.Q 7.52e-19
C13374 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_891_329# -3.3e-20
C13375 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# -0.00106f
C13376 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# -3.79e-20
C13377 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# -4.66e-20
C13378 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__inv_1_32/Y 2.47e-20
C13379 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# V_LOW 0.00727f
C13380 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_28/Y 0.0316f
C13381 sky130_fd_sc_hd__inv_1_64/A CLOCK_GEN.SR_Op.Q 0.017f
C13382 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 6.82e-20
C13383 sky130_fd_sc_hd__inv_16_26/A sky130_fd_sc_hd__inv_16_7/Y 0.0487f
C13384 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 6.27e-19
C13385 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# sky130_fd_sc_hd__inv_1_40/Y 9.3e-22
C13386 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 0.028f
C13387 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_1_1/Y 3.02e-20
C13388 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF2.Q 5.17e-20
C13389 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# -0.00592f
C13390 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 6.94e-19
C13391 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 0.00803f
C13392 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00116f
C13393 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 5.52e-19
C13394 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_557_413# 4.54e-19
C13395 sky130_fd_sc_hd__inv_1_24/Y V_LOW 0.23f
C13396 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_16_4/Y 0.00897f
C13397 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00379f
C13398 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__inv_1_50/Y 6.02e-19
C13399 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 1.46e-20
C13400 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_0/HI 0.0266f
C13401 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__conb_1_39/LO 9.91e-20
C13402 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__inv_16_41/Y 0.0299f
C13403 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_1_19/A 5.5e-20
C13404 sky130_fd_sc_hd__dfbbn_1_37/Q_N V_LOW -0.00245f
C13405 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_1_36/Y 2.89e-21
C13406 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# V_LOW -0.103f
C13407 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__conb_1_31/HI 1.96e-21
C13408 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# 8.66e-21
C13409 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.00576f
C13410 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# V_LOW -6.55e-19
C13411 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# V_LOW -0.00266f
C13412 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 9.9e-21
C13413 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# -1.44e-20
C13414 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 4.54e-20
C13415 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_59/Y 2.65e-21
C13416 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# V_LOW 2.26e-20
C13417 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__inv_1_30/Y 3.7e-20
C13418 RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 3.97e-19
C13419 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_27/LO 2.7e-19
C13420 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# -2.52e-19
C13421 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -0.0114f
C13422 sky130_fd_sc_hd__conb_1_23/LO FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0431f
C13423 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__inv_1_60/Y 2e-19
C13424 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__conb_1_28/HI 2.2e-19
C13425 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__conb_1_4/LO 2.15e-19
C13426 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# Reset 0.00165f
C13427 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_11/LO 3.51e-20
C13428 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_41/HI 0.45f
C13429 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_1_44/A 0.00123f
C13430 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# 0.00147f
C13431 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 7.52e-21
C13432 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# V_LOW 3.56e-20
C13433 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# V_LOW 0.0114f
C13434 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 5.1e-20
C13435 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 8.37e-20
C13436 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0415f
C13437 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__nor2_1_0/Y 0.00287f
C13438 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__inv_16_40/Y 4.07e-20
C13439 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_38/LO 4.79e-19
C13440 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.23e-19
C13441 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 8.97e-20
C13442 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 7.39e-20
C13443 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 8.97e-20
C13444 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0.0127f
C13445 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 7.39e-20
C13446 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 0.0452f
C13447 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_50/HI 0.171f
C13448 FALLING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 1.44f
C13449 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.00106f
C13450 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 5.05e-19
C13451 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00122f
C13452 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 4.66e-19
C13453 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 7.6e-21
C13454 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.18e-22
C13455 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_1_43/Y 3.28e-20
C13456 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 6.87e-19
C13457 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_12/LO 3.56e-21
C13458 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 6.39e-19
C13459 FULL_COUNTER.COUNT_SUB_DFF2.Q Reset 1.97f
C13460 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 5.65e-19
C13461 sky130_fd_sc_hd__nand2_8_4/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 6.04e-20
C13462 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 2.02e-19
C13463 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0163f
C13464 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_16_42/Y 0.0164f
C13465 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_16_40/Y 2.93e-22
C13466 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# -1.24e-20
C13467 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_31/HI 9.47e-21
C13468 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# V_LOW 2.26e-20
C13469 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 5.68e-20
C13470 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 1.08e-20
C13471 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_1_8/Y 0.00345f
C13472 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 7.24e-19
C13473 sky130_fd_sc_hd__dfbbn_1_15/Q_N FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00669f
C13474 sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__inv_1_26/Y 2.5e-21
C13475 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 0.637f
C13476 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_3/HI 1.61e-19
C13477 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 8.92e-21
C13478 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_22/A 0.068f
C13479 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00127f
C13480 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 8.31e-19
C13481 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 8.68e-20
C13482 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 7.27e-19
C13483 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_45/a_381_47# 2.28e-19
C13484 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_1_2/Y 0.0317f
C13485 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# -0.00592f
C13486 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0216f
C13487 sky130_fd_sc_hd__conb_1_36/LO Reset 2.44e-19
C13488 sky130_fd_sc_hd__inv_1_27/Y V_LOW 0.463f
C13489 sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# sky130_fd_sc_hd__inv_1_28/Y 1.57e-19
C13490 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# V_LOW 2.27e-19
C13491 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 9.58e-21
C13492 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_64/A 0.00106f
C13493 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00777f
C13494 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00498f
C13495 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 8e-21
C13496 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# V_LOW 0.00224f
C13497 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_791_47# 9.26e-20
C13498 sky130_fd_sc_hd__inv_1_61/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0117f
C13499 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/Q_N -6.48e-19
C13500 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 3.35e-19
C13501 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__conb_1_17/HI 0.0021f
C13502 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 0.0149f
C13503 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 3.27e-19
C13504 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__inv_1_30/Y 0.0146f
C13505 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__inv_1_50/Y 0.00308f
C13506 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_891_329# 1.5e-21
C13507 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_19/A 0.0101f
C13508 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# -4.66e-20
C13509 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# -3.79e-20
C13510 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# -0.0128f
C13511 sky130_fd_sc_hd__dfbbn_1_44/a_581_47# sky130_fd_sc_hd__inv_16_41/Y 0.00167f
C13512 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.76e-19
C13513 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nand2_8_9/A 6.43e-20
C13514 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# V_LOW -2.68e-19
C13515 sky130_fd_sc_hd__inv_1_41/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0911f
C13516 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__inv_1_32/Y 3.42e-20
C13517 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_35/Y 0.00465f
C13518 sky130_fd_sc_hd__nand3_1_2/Y CLOCK_GEN.SR_Op.Q 0.173f
C13519 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_36/Y 1.48e-20
C13520 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.002f
C13521 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# sky130_fd_sc_hd__inv_1_35/Y 3.72e-20
C13522 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 4.35e-19
C13523 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00608f
C13524 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# V_LOW 0.00124f
C13525 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00111f
C13526 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_51/Y 6.79e-20
C13527 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.57e-19
C13528 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# -1.76e-19
C13529 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# -6.29e-19
C13530 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_891_329# -2.46e-19
C13531 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_557_413# -3.67e-20
C13532 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__inv_1_44/A 7.36e-21
C13533 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_2_0/A 0.0422f
C13534 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_8/HI 0.0242f
C13535 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 7.04e-19
C13536 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 4.85e-21
C13537 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0.00147f
C13538 sky130_fd_sc_hd__nand2_8_8/A sky130_fd_sc_hd__nand2_1_5/Y 5.46e-20
C13539 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__inv_1_60/Y 0.0977f
C13540 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# sky130_fd_sc_hd__nor2_1_0/Y 4.49e-21
C13541 sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 2.11e-20
C13542 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__inv_1_2/Y 3.91e-20
C13543 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.01e-19
C13544 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# -4.66e-20
C13545 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_381_47# -3.79e-20
C13546 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_34/HI 0.0147f
C13547 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 4.17e-20
C13548 sky130_fd_sc_hd__conb_1_16/HI FULL_COUNTER.COUNT_SUB_DFF14.Q 0.841f
C13549 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_1_29/Y 3.53e-20
C13550 FALLING_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0314f
C13551 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 8.81e-20
C13552 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00604f
C13553 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 5.91e-20
C13554 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_581_47# -2.6e-20
C13555 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 5.91e-19
C13556 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 1.34e-20
C13557 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# sky130_fd_sc_hd__inv_1_8/Y 2.02e-19
C13558 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00196f
C13559 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0.00196f
C13560 sky130_fd_sc_hd__conb_1_30/HI RISING_COUNTER.COUNT_SUB_DFF10.Q 0.106f
C13561 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_49/A 7.23e-19
C13562 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0293f
C13563 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00103f
C13564 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# V_LOW 4.8e-20
C13565 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# 5.94e-19
C13566 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.0381f
C13567 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 2.58e-19
C13568 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_42/LO 9.95e-20
C13569 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__inv_1_32/Y 3.68e-21
C13570 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_58/Y 0.00293f
C13571 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__conb_1_34/LO 2.77e-20
C13572 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# V_LOW 1.79e-20
C13573 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 0.0149f
C13574 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_1_1/Y 5.49e-19
C13575 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__inv_1_62/Y 0.195f
C13576 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_48/Y 8.2e-21
C13577 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_557_413# -0.0012f
C13578 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# -0.0309f
C13579 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 0.199f
C13580 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# V_LOW -0.00389f
C13581 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00125f
C13582 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__conb_1_47/HI 0.00139f
C13583 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.69e-21
C13584 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 8.47e-19
C13585 sky130_fd_sc_hd__inv_1_35/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.17e-19
C13586 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__conb_1_17/HI 8.64e-21
C13587 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.18e-20
C13588 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# sky130_fd_sc_hd__inv_1_35/Y 1.44e-21
C13589 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__nand3_1_2/Y 1.45e-20
C13590 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_66/Y 6.56e-22
C13591 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__conb_1_12/HI 0.00353f
C13592 sky130_fd_sc_hd__inv_1_3/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00117f
C13593 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# V_LOW 6.75e-19
C13594 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.00581f
C13595 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# -1.69e-19
C13596 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00116f
C13597 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_2_0/A 0.0448f
C13598 sky130_fd_sc_hd__conb_1_50/LO FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0173f
C13599 sky130_fd_sc_hd__inv_1_67/A sky130_fd_sc_hd__inv_1_66/A 0.408f
C13600 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_44/A 0.143f
C13601 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_27/Y 0.00204f
C13602 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__inv_1_41/Y 0.00931f
C13603 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_5/HI 1.07e-21
C13604 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__conb_1_24/HI 9.41e-22
C13605 sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__inv_1_24/Y 2.17e-19
C13606 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# -1.27e-19
C13607 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_66/A 1.2e-19
C13608 sky130_fd_sc_hd__nand2_1_3/Y V_LOW -0.00556f
C13609 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_17/HI 0.0251f
C13610 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__conb_1_38/HI 0.00399f
C13611 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00469f
C13612 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00227f
C13613 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__conb_1_27/HI 0.0185f
C13614 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_16_42/Y 1.61e-19
C13615 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__conb_1_20/HI 0.0037f
C13616 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_941_21# 7.38e-19
C13617 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_1_43/Y 2.99e-21
C13618 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_891_329# 5.62e-21
C13619 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00155f
C13620 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# -0.00409f
C13621 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# -0.0103f
C13622 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0397f
C13623 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.03e-20
C13624 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 0.0234f
C13625 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__inv_1_21/Y 4.18e-19
C13626 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 3.88e-19
C13627 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 4.12e-19
C13628 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 5.94e-19
C13629 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.88e-19
C13630 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_29/Y 7.41e-20
C13631 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00158f
C13632 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_34/LO 0.00185f
C13633 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# sky130_fd_sc_hd__conb_1_21/HI 0.00107f
C13634 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# sky130_fd_sc_hd__inv_1_31/Y 2.03e-21
C13635 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.201f
C13636 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0.00171f
C13637 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__conb_1_24/HI -0.00907f
C13638 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__conb_1_17/LO 3.38e-20
C13639 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_38/HI 0.0887f
C13640 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__inv_1_38/Y 0.0101f
C13641 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__inv_1_58/Y 0.0141f
C13642 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__conb_1_16/HI 8.19e-22
C13643 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_3/LO 0.00131f
C13644 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# V_LOW 0.00244f
C13645 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 6.94e-19
C13646 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.00116f
C13647 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 0.00803f
C13648 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 5.52e-19
C13649 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# -4.36e-19
C13650 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_2_0/A 2.28e-20
C13651 V_HIGH FULL_COUNTER.COUNT_SUB_DFF0.Q 1.33f
C13652 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.93e-20
C13653 sky130_fd_sc_hd__inv_16_6/A FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.121f
C13654 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_46/A 7.14e-19
C13655 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__inv_1_33/Y 1.56e-20
C13656 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0132f
C13657 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 5.88e-21
C13658 sky130_fd_sc_hd__conb_1_11/LO FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00344f
C13659 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.35e-19
C13660 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__conb_1_12/HI 0.0045f
C13661 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.00911f
C13662 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_581_47# -7.91e-19
C13663 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# V_LOW 2.94e-20
C13664 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__conb_1_4/HI 0.00169f
C13665 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0126f
C13666 sky130_fd_sc_hd__dfbbn_1_24/Q_N FALLING_COUNTER.COUNT_SUB_DFF15.Q 0.0338f
C13667 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 1.59e-19
C13668 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0.00637f
C13669 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 3.03e-21
C13670 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 8.98e-19
C13671 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 6.89e-19
C13672 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__conb_1_5/HI 2.42e-21
C13673 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_49/Y 0.377f
C13674 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.00141f
C13675 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -6.23e-21
C13676 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -1.42e-32
C13677 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_381_47# -0.00393f
C13678 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_581_47# -2.6e-20
C13679 sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF14.Q 9.9e-19
C13680 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__inv_1_66/A 3.86e-20
C13681 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# V_LOW 3.56e-20
C13682 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_2/Q_N -1.42e-32
C13683 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__conb_1_17/HI 7.82e-19
C13684 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0.0107f
C13685 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 0.00182f
C13686 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 2.69e-19
C13687 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 1.7e-20
C13688 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 4.64e-19
C13689 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__inv_1_25/Y 9.58e-19
C13690 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# sky130_fd_sc_hd__conb_1_20/HI 2.78e-21
C13691 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# sky130_fd_sc_hd__conb_1_27/HI -0.00263f
C13692 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__conb_1_46/HI 4.84e-20
C13693 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__inv_1_45/Y 7.41e-22
C13694 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 1.96e-19
C13695 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# V_LOW 1.38e-19
C13696 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__conb_1_37/HI 8.76e-20
C13697 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 3.87e-20
C13698 sky130_fd_sc_hd__inv_1_22/Y Reset 0.036f
C13699 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# -0.00235f
C13700 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# -7.93e-19
C13701 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_33/Y 0.0366f
C13702 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_50/HI 7.92e-21
C13703 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# -5.14e-19
C13704 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__inv_1_7/Y 5.71e-19
C13705 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00477f
C13706 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.56e-21
C13707 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 7.09e-20
C13708 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__inv_1_34/Y 0.00575f
C13709 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 1.03e-20
C13710 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 4.97e-20
C13711 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_26/Y 0.0602f
C13712 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 2.24e-20
C13713 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__inv_1_29/Y 5.18e-20
C13714 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# V_LOW 2.26e-20
C13715 FULL_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF8.Q 1.3e-19
C13716 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.49f
C13717 RISING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.26e-19
C13718 sky130_fd_sc_hd__inv_1_52/A Reset 7.14e-19
C13719 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 0.329f
C13720 sky130_fd_sc_hd__inv_16_42/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0963f
C13721 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_1_2/A 0.195f
C13722 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF9.Q 1.51e-20
C13723 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_8_0/Y 2.07e-20
C13724 sky130_fd_sc_hd__conb_1_49/LO FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00968f
C13725 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.03e-19
C13726 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.87e-21
C13727 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_1_10/Y 1.6e-19
C13728 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__conb_1_51/HI 3.34e-20
C13729 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__conb_1_12/HI -0.0614f
C13730 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__conb_1_5/HI 1.83e-20
C13731 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__conb_1_24/HI -9.71e-19
C13732 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 0.002f
C13733 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# sky130_fd_sc_hd__inv_1_38/Y 7.18e-21
C13734 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00137f
C13735 sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF14.Q 0.149f
C13736 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 2.43e-20
C13737 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_47/Y 7.92e-20
C13738 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00116f
C13739 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_647_21# -0.00155f
C13740 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_473_413# -0.00536f
C13741 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_26/LO 2.42e-21
C13742 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# V_LOW 2.94e-20
C13743 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_10/HI 2.38e-19
C13744 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# 3.35e-19
C13745 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 6.28e-20
C13746 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.0029f
C13747 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 0.00106f
C13748 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 0.0035f
C13749 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_29/HI 0.109f
C13750 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00421f
C13751 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 3.77e-19
C13752 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 6.78e-19
C13753 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__conb_1_51/HI 2.73e-20
C13754 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1_66/A 3.36e-20
C13755 sky130_fd_sc_hd__inv_16_7/A sky130_fd_sc_hd__inv_16_8/A 0.0121f
C13756 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_16_40/Y 0.00162f
C13757 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 0.001f
C13758 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_33/Y 0.136f
C13759 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__conb_1_44/HI 0.00314f
C13760 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 7.18e-19
C13761 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__conb_1_43/HI 0.0243f
C13762 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# Reset 0.00653f
C13763 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# -0.00149f
C13764 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# -0.00441f
C13765 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 8e-21
C13766 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00224f
C13767 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 7.09e-19
C13768 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 3.67e-21
C13769 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# -1.64e-20
C13770 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__conb_1_12/HI 0.0028f
C13771 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_28/Y 2.64e-19
C13772 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__conb_1_4/HI 1.17e-19
C13773 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0257f
C13774 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_24/Y 0.00558f
C13775 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 5.28e-19
C13776 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 2.06e-19
C13777 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 7.01e-19
C13778 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 7.04e-19
C13779 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# -5.54e-21
C13780 sky130_fd_sc_hd__conb_1_51/LO V_LOW 0.0459f
C13781 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.36e-19
C13782 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 6.13e-20
C13783 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_16_42/Y 0.0227f
C13784 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00344f
C13785 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0891f
C13786 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# 3.57e-20
C13787 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0063f
C13788 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_1_12/Y 2.89e-21
C13789 sky130_fd_sc_hd__conb_1_40/LO V_LOW 0.0881f
C13790 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -1.03e-19
C13791 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# -3.86e-20
C13792 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# V_LOW 0.0109f
C13793 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__inv_16_41/Y 1.53e-20
C13794 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 0.0446f
C13795 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# V_LOW 2.26e-20
C13796 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__conb_1_46/HI 9.36e-20
C13797 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_18/HI 2.4e-19
C13798 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# V_LOW -0.006f
C13799 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/Q_N -4.24e-20
C13800 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__conb_1_5/HI 2.59e-20
C13801 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# -1.76e-19
C13802 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_381_47# 1.22e-20
C13803 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__inv_1_12/Y 9.63e-19
C13804 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 2.36e-21
C13805 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00111f
C13806 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# -0.00336f
C13807 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# -3.79e-20
C13808 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 9.89e-21
C13809 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF6.Q -5.45e-20
C13810 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# sky130_fd_sc_hd__conb_1_11/HI 0.00519f
C13811 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 2.47e-19
C13812 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 7.33e-19
C13813 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# V_LOW -0.00266f
C13814 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.88e-19
C13815 sky130_fd_sc_hd__inv_1_46/A Reset 4.6e-19
C13816 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF2.Q 1.19e-20
C13817 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_1_7/Y 0.0017f
C13818 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 2.93e-21
C13819 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 3.94e-19
C13820 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.48e-19
C13821 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 2.95e-22
C13822 sky130_fd_sc_hd__inv_1_66/Y CLOCK_GEN.SR_Op.Q 0.0239f
C13823 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 2.27e-20
C13824 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00157f
C13825 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__conb_1_24/HI 4.59e-21
C13826 V_SENSE sky130_fd_sc_hd__inv_16_49/A 0.799f
C13827 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.119f
C13828 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# sky130_fd_sc_hd__inv_1_37/Y 0.00135f
C13829 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.88e-19
C13830 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.83e-19
C13831 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_51/Y 4.23e-21
C13832 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__conb_1_32/HI 0.00249f
C13833 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 7.06e-19
C13834 sky130_fd_sc_hd__conb_1_16/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 0.176f
C13835 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 3.58e-19
C13836 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.00996f
C13837 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# V_LOW 0.0659f
C13838 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_10/HI -4.84e-20
C13839 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.53e-21
C13840 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.55e-19
C13841 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 5.74e-20
C13842 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 0.00104f
C13843 FALLING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0485f
C13844 sky130_fd_sc_hd__conb_1_35/HI CLOCK_GEN.SR_Op.Q 9.98e-20
C13845 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0.0274f
C13846 sky130_fd_sc_hd__dfbbn_1_49/Q_N FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.27e-19
C13847 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_38/HI 4.09e-22
C13848 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__inv_1_50/Y 1.07e-20
C13849 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 3.57e-20
C13850 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 2.82e-21
C13851 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 8.83e-19
C13852 sky130_fd_sc_hd__conb_1_26/LO V_LOW 0.0718f
C13853 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# -9.62e-19
C13854 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_48/A 8.88e-19
C13855 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# 0.00477f
C13856 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# sky130_fd_sc_hd__conb_1_44/HI -1.17e-19
C13857 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.38e-19
C13858 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# 6.49e-19
C13859 sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_16_19/Y 0.00907f
C13860 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# Reset 0.00472f
C13861 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0364f
C13862 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# -0.00141f
C13863 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00425f
C13864 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# CLOCK_GEN.SR_Op.Q 7.54e-20
C13865 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 0.0015f
C13866 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__conb_1_37/HI 0.00391f
C13867 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# sky130_fd_sc_hd__conb_1_37/HI -6.57e-19
C13868 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# sky130_fd_sc_hd__inv_16_42/Y 2.39e-20
C13869 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.41e-21
C13870 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_44/A 0.132f
C13871 sky130_fd_sc_hd__conb_1_37/LO V_LOW 0.125f
C13872 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.036f
C13873 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 8.8e-22
C13874 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 2.14e-20
C13875 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.36e-19
C13876 RISING_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0241f
C13877 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -0.00907f
C13878 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00293f
C13879 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 0.00225f
C13880 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 4.33e-19
C13881 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_1_30/Y 0.0248f
C13882 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_38/HI 0.273f
C13883 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 1.96e-20
C13884 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.273f
C13885 RISING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0187f
C13886 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 1.2e-19
C13887 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__inv_16_40/Y 0.0311f
C13888 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__inv_1_36/Y 0.00977f
C13889 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_10/Y 0.023f
C13890 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 0.0148f
C13891 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# -2.53e-20
C13892 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_44/A 1.44e-20
C13893 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.95e-19
C13894 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_46/LO 1.37e-20
C13895 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_47/Y 0.222f
C13896 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_39/Y 0.0367f
C13897 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# -2.57e-20
C13898 sky130_fd_sc_hd__inv_1_47/A FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0676f
C13899 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__inv_16_41/Y 3.52e-21
C13900 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_473_413# -0.00591f
C13901 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_647_21# -6.43e-20
C13902 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# sky130_fd_sc_hd__conb_1_46/HI 2.47e-19
C13903 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__conb_1_18/HI 2.62e-20
C13904 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00146f
C13905 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# V_LOW 2.94e-20
C13906 FALLING_COUNTER.COUNT_SUB_DFF11.Q V_LOW 2.06f
C13907 sky130_fd_sc_hd__inv_1_35/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 7.73e-20
C13908 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 0.00138f
C13909 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_40/Y 0.00231f
C13910 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 9.31e-20
C13911 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# 1.35e-19
C13912 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__conb_1_21/HI 0.0122f
C13913 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_22/Y 0.00305f
C13914 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 1.07e-19
C13915 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# -0.00138f
C13916 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -2.18e-19
C13917 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -5.54e-21
C13918 sky130_fd_sc_hd__inv_1_24/A Reset 4.83e-19
C13919 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 6.46e-24
C13920 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_39/HI 1.9e-20
C13921 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# V_LOW 4.8e-20
C13922 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00626f
C13923 sky130_fd_sc_hd__inv_1_3/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0246f
C13924 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_44/A 0.0242f
C13925 sky130_fd_sc_hd__conb_1_29/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00105f
C13926 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_1_49/Y 0.00623f
C13927 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_32/HI 0.00218f
C13928 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_5/HI -5.52e-19
C13929 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__conb_1_7/HI 9.67e-20
C13930 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__inv_16_40/Y 2.62e-19
C13931 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__conb_1_24/HI 4.28e-21
C13932 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.03e-21
C13933 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__conb_1_46/HI 1.05e-20
C13934 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__conb_1_19/HI 1.92e-20
C13935 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__inv_1_44/A 0.0227f
C13936 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0356f
C13937 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_55/Y 0.227f
C13938 sky130_fd_sc_hd__dfbbn_1_28/a_581_47# sky130_fd_sc_hd__conb_1_32/HI 2.13e-19
C13939 sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__dfbbn_1_10/a_791_47# -0.01f
C13940 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 0.00971f
C13941 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__conb_1_12/HI 3.27e-21
C13942 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 2.38e-20
C13943 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 7.44e-21
C13944 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 4.58e-19
C13945 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# V_LOW 2.94e-20
C13946 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_891_329# -2.2e-20
C13947 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# -0.00953f
C13948 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__conb_1_25/HI 0.00535f
C13949 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 3.97e-23
C13950 sky130_fd_sc_hd__inv_1_42/Y V_LOW 0.0469f
C13951 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_1_13/Y 0.00698f
C13952 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__conb_1_23/HI 0.00211f
C13953 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_31/Y 0.261f
C13954 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0.00127f
C13955 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 8.32e-19
C13956 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_35/HI 1.05e-20
C13957 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_45/A 0.136f
C13958 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_21/HI 0.0184f
C13959 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 6.38e-20
C13960 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 1.54e-19
C13961 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 5.26e-21
C13962 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# V_LOW 0.0122f
C13963 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# -9.32e-20
C13964 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_10/Y 0.00274f
C13965 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# V_LOW 1.38e-19
C13966 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0241f
C13967 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_48/HI 4.18e-21
C13968 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 0.00725f
C13969 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 0.0714f
C13970 sky130_fd_sc_hd__inv_1_52/Y CLOCK_GEN.SR_Op.Q 4.68e-19
C13971 sky130_fd_sc_hd__inv_16_40/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0697f
C13972 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__nand2_8_4/Y 1.01e-21
C13973 sky130_fd_sc_hd__dfbbn_1_32/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00216f
C13974 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/Q_N -9.56e-20
C13975 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# V_LOW 0.00126f
C13976 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# CLOCK_GEN.SR_Op.Q 1.49e-20
C13977 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 9.44e-19
C13978 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 6.21e-20
C13979 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0472f
C13980 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 2.05e-19
C13981 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 5.45e-19
C13982 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/Q_N -4.78e-20
C13983 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q -3.39e-20
C13984 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# 1.55e-20
C13985 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 6.25e-19
C13986 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# -9.71e-19
C13987 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.00211f
C13988 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# V_LOW 0.0154f
C13989 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__inv_1_40/Y 0.025f
C13990 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__conb_1_33/HI -0.00106f
C13991 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 3.72e-19
C13992 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__inv_16_40/Y 0.00415f
C13993 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 4.98e-20
C13994 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__conb_1_9/HI 6.19e-20
C13995 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_56/Y 0.0768f
C13996 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_44/A 0.00242f
C13997 sky130_fd_sc_hd__inv_4_0/A FULL_COUNTER.COUNT_SUB_DFF0.Q 2.81e-21
C13998 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00218f
C13999 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 0.00521f
C14000 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# -1.44e-20
C14001 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 0.00265f
C14002 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# -0.0266f
C14003 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_557_413# -0.0012f
C14004 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 2.85e-19
C14005 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__conb_1_31/HI -0.00201f
C14006 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__inv_1_69/Y 0.00481f
C14007 sky130_fd_sc_hd__conb_1_26/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 0.002f
C14008 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 4.15e-19
C14009 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__conb_1_18/HI 7.43e-21
C14010 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.84e-19
C14011 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# V_LOW 0.0257f
C14012 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# sky130_fd_sc_hd__inv_1_40/Y 1.57e-21
C14013 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00212f
C14014 sky130_fd_sc_hd__conb_1_35/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0209f
C14015 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__conb_1_5/HI 1.01e-19
C14016 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# sky130_fd_sc_hd__conb_1_28/HI 0.00135f
C14017 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__inv_1_29/Y 7.36e-19
C14018 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# -9.32e-20
C14019 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_1_25/Y 2.26e-20
C14020 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_647_21# 0.0238f
C14021 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_26/Y 0.0248f
C14022 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__conb_1_5/HI -0.0127f
C14023 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_1_61/Y 1.3e-19
C14024 sky130_fd_sc_hd__nand2_8_9/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 3.63e-19
C14025 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 6.03e-19
C14026 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.78e-19
C14027 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.32e-19
C14028 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0262f
C14029 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/Q_N 7.16e-21
C14030 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_1_2/Y 5.3e-19
C14031 sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 1.27e-20
C14032 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__inv_1_44/A 0.00397f
C14033 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_23/HI 0.00301f
C14034 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__conb_1_19/LO 0.00434f
C14035 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__inv_1_13/Y 7.45e-21
C14036 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00787f
C14037 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 2.37e-20
C14038 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# -0.0129f
C14039 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# -0.00864f
C14040 FALLING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 7.51e-19
C14041 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# 2.65e-19
C14042 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# -0.055f
C14043 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__nand2_1_2/A 3.88e-19
C14044 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# -0.00592f
C14045 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__conb_1_25/HI 0.0191f
C14046 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.341f
C14047 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# sky130_fd_sc_hd__inv_1_13/Y 4.05e-19
C14048 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_1_39/Y 9.87e-20
C14049 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 1.8e-20
C14050 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__conb_1_8/LO 2.45e-20
C14051 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__dfbbn_1_13/a_557_413# 4.43e-19
C14052 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# sky130_fd_sc_hd__inv_1_33/Y 4.1e-21
C14053 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_1_66/A 3.05e-20
C14054 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_31/Y 0.147f
C14055 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__inv_1_50/Y 5.85e-22
C14056 sky130_fd_sc_hd__inv_16_55/A sky130_fd_sc_hd__inv_16_50/A 8.88e-19
C14057 sky130_fd_sc_hd__inv_16_15/A V_LOW 0.241f
C14058 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_4_0/A 4.63e-19
C14059 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/Q_N -4.78e-20
C14060 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__conb_1_45/HI -4.99e-19
C14061 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_16/LO 0.00195f
C14062 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# sky130_fd_sc_hd__inv_1_10/Y 7.48e-20
C14063 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00411f
C14064 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__conb_1_48/HI 2.14e-20
C14065 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF14.Q 5.54e-19
C14066 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# 4.91e-20
C14067 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# 2.85e-19
C14068 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_36/LO 6.66e-19
C14069 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 0.005f
C14070 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 1.29e-20
C14071 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# V_LOW -1.39e-35
C14072 FULL_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 1.61e-20
C14073 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 0.119f
C14074 FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00139f
C14075 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 4.85e-21
C14076 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 2.78e-20
C14077 RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.155f
C14078 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_16_4/Y 2.26e-21
C14079 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0238f
C14080 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 4.21e-19
C14081 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_52/A 2.22e-19
C14082 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00768f
C14083 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_10/Y 0.38f
C14084 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__conb_1_6/HI 1.22e-20
C14085 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_42/Q_N -2.17e-19
C14086 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# V_LOW 2.26e-20
C14087 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0211f
C14088 sky130_fd_sc_hd__conb_1_40/HI V_LOW 0.0432f
C14089 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# -1.62e-20
C14090 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# -2.37e-19
C14091 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# V_LOW 1.79e-20
C14092 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_41/a_381_47# 0.00315f
C14093 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__conb_1_33/HI -2.07e-19
C14094 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__dfbbn_1_15/Q_N 1.16e-19
C14095 sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 0.106f
C14096 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.91e-19
C14097 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_7/HI 5.27e-21
C14098 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_22/a_791_47# 4.19e-20
C14099 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# -5.42e-19
C14100 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# sky130_fd_sc_hd__conb_1_31/HI -7.2e-19
C14101 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0298f
C14102 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_1_41/Y 1.37e-19
C14103 sky130_fd_sc_hd__conb_1_36/LO FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00312f
C14104 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8e-20
C14105 sky130_fd_sc_hd__dfbbn_1_50/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00126f
C14106 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_45/Y 3.87e-20
C14107 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.09e-19
C14108 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_7/LO 1e-19
C14109 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# V_LOW 3.84e-19
C14110 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.72e-19
C14111 sky130_fd_sc_hd__nand3_1_2/a_193_47# CLOCK_GEN.SR_Op.Q 2.34e-19
C14112 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_891_329# -2.2e-20
C14113 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# -4.72e-19
C14114 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__inv_1_39/Y 4.18e-20
C14115 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/Q_N -4.78e-20
C14116 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_16/HI 5.53e-19
C14117 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0174f
C14118 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_38/a_581_47# 0.00101f
C14119 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00211f
C14120 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF14.Q 8.77e-19
C14121 RISING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.68f
C14122 sky130_fd_sc_hd__inv_16_32/Y sky130_fd_sc_hd__inv_16_28/Y 0.153f
C14123 sky130_fd_sc_hd__inv_16_15/A sky130_fd_sc_hd__inv_16_9/Y 0.00211f
C14124 sky130_fd_sc_hd__conb_1_13/HI FULL_COUNTER.COUNT_SUB_DFF18.Q 0.196f
C14125 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__conb_1_11/LO 0.0656f
C14126 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_32/Y 1.08e-20
C14127 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__conb_1_2/HI 0.00147f
C14128 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00277f
C14129 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.0106f
C14130 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 1.34e-19
C14131 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 0.023f
C14132 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 1.1e-19
C14133 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.21e-20
C14134 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__inv_1_2/Y 0.00306f
C14135 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__conb_1_19/HI 1.68e-20
C14136 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# V_LOW 0.0115f
C14137 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 9.02e-20
C14138 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# Reset 0.00286f
C14139 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_40/Y 0.127f
C14140 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# sky130_fd_sc_hd__conb_1_23/HI 5.75e-19
C14141 sky130_fd_sc_hd__conb_1_27/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 1.46e-19
C14142 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_9/A 2.58e-20
C14143 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.00124f
C14144 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__conb_1_45/LO 0.00221f
C14145 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0131f
C14146 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__inv_1_1/Y 0.00163f
C14147 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 9.72e-20
C14148 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 2.13e-19
C14149 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 1.77e-19
C14150 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__inv_1_60/Y 0.00975f
C14151 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# -0.0162f
C14152 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__conb_1_30/HI 9.79e-19
C14153 sky130_fd_sc_hd__conb_1_23/HI V_LOW 0.221f
C14154 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 3.23e-20
C14155 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_1_39/Y 5.82e-20
C14156 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# V_LOW 0.0203f
C14157 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__inv_1_14/Y 0.00318f
C14158 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_48/Y 1.71e-19
C14159 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__conb_1_41/HI 0.00164f
C14160 sky130_fd_sc_hd__dfbbn_1_10/Q_N FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00155f
C14161 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_22/A 2.57e-19
C14162 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 8.81e-20
C14163 sky130_fd_sc_hd__inv_16_14/Y V_LOW 0.316f
C14164 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 3.61e-21
C14165 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.81e-20
C14166 sky130_fd_sc_hd__dfbbn_1_1/Q_N V_LOW -0.00509f
C14167 RISING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.05e-20
C14168 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 8.17e-19
C14169 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_21/Y 5.14e-19
C14170 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 2.65e-20
C14171 sky130_fd_sc_hd__inv_1_32/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.769f
C14172 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00378f
C14173 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__inv_1_10/Y 0.00186f
C14174 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__conb_1_50/HI 1.68e-19
C14175 sky130_fd_sc_hd__nand2_8_9/A sky130_fd_sc_hd__inv_1_66/A 0.0347f
C14176 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# sky130_fd_sc_hd__conb_1_6/HI 1.35e-19
C14177 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 3.11e-19
C14178 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 0.0063f
C14179 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 0.00902f
C14180 sky130_fd_sc_hd__inv_16_32/A sky130_fd_sc_hd__inv_16_28/Y 7.06e-19
C14181 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# -1.66e-19
C14182 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 0.0182f
C14183 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_53/Y 8.73e-21
C14184 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__inv_1_28/Y 3.69e-19
C14185 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__inv_2_0/A 0.00292f
C14186 sky130_fd_sc_hd__inv_16_49/A CLOCK_GEN.SR_Op.Q 0.0271f
C14187 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__conb_1_31/HI 5.56e-19
C14188 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__inv_1_41/Y 4.93e-20
C14189 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__inv_1_21/Y 1.56e-19
C14190 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_66/A 2.01e-20
C14191 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# -2.66e-19
C14192 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# -2.52e-19
C14193 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__conb_1_39/HI 0.00275f
C14194 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# 1.42e-32
C14195 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# -0.00471f
C14196 sky130_fd_sc_hd__conb_1_30/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 2.11e-19
C14197 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_473_413# -0.00458f
C14198 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_647_21# -0.00431f
C14199 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.06e-20
C14200 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_55/Y 0.267f
C14201 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 7.13e-22
C14202 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 6.54e-20
C14203 V_SENSE sky130_fd_sc_hd__inv_16_6/Y 0.0168f
C14204 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_66/A 0.21f
C14205 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_67/A 1.37e-20
C14206 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__conb_1_2/HI 5.05e-19
C14207 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# V_LOW 4.8e-20
C14208 sky130_fd_sc_hd__inv_16_8/Y V_LOW 0.242f
C14209 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 2.66e-19
C14210 sky130_fd_sc_hd__inv_16_14/Y sky130_fd_sc_hd__inv_16_9/Y 1.28e-19
C14211 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 0.00496f
C14212 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 1.48e-20
C14213 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.34e-20
C14214 sky130_fd_sc_hd__inv_1_36/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 1.27e-20
C14215 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# V_LOW -3.78e-19
C14216 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.5e-21
C14217 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# V_LOW -0.0176f
C14218 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# V_LOW 2.26e-20
C14219 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 0.00232f
C14220 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# -0.0672f
C14221 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00124f
C14222 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# V_LOW 0.0323f
C14223 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__conb_1_45/LO 1.75e-19
C14224 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00102f
C14225 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00292f
C14226 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.68e-19
C14227 sky130_fd_sc_hd__conb_1_19/LO V_LOW 0.0962f
C14228 sky130_fd_sc_hd__inv_1_47/A FULL_COUNTER.COUNT_SUB_DFF0.Q 2.27e-19
C14229 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__conb_1_9/HI 1.93e-19
C14230 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# sky130_fd_sc_hd__inv_1_60/Y 2.05e-21
C14231 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__dfbbn_1_38/a_473_413# 3.38e-20
C14232 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# sky130_fd_sc_hd__inv_16_41/Y 1.01e-19
C14233 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# V_LOW -0.309f
C14234 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__inv_1_39/Y 0.00538f
C14235 V_SENSE sky130_fd_sc_hd__inv_16_33/Y 0.00177f
C14236 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# V_LOW 2.94e-20
C14237 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# sky130_fd_sc_hd__inv_1_14/Y 1.07e-21
C14238 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__inv_1_8/Y 8.34e-20
C14239 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 0.0199f
C14240 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 0.00721f
C14241 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# 7.12e-19
C14242 sky130_fd_sc_hd__dfbbn_1_46/a_581_47# sky130_fd_sc_hd__conb_1_41/HI 2.47e-19
C14243 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_0/Y 0.038f
C14244 Reset FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.193f
C14245 sky130_fd_sc_hd__nand2_8_4/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0303f
C14246 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_45/Q_N 0.00178f
C14247 sky130_fd_sc_hd__inv_1_3/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0278f
C14248 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.47e-19
C14249 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_47/Y 5.67e-20
C14250 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_1_61/Y 5.29e-20
C14251 sky130_fd_sc_hd__conb_1_29/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00162f
C14252 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# sky130_fd_sc_hd__conb_1_4/HI 4.06e-19
C14253 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 9.34e-19
C14254 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# sky130_fd_sc_hd__inv_1_38/Y 0.00119f
C14255 sky130_fd_sc_hd__dfbbn_1_30/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00424f
C14256 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__conb_1_26/HI 0.0213f
C14257 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# -4.66e-20
C14258 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# -3.79e-20
C14259 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__conb_1_16/LO 1.03e-20
C14260 sky130_fd_sc_hd__inv_1_69/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 8.34e-19
C14261 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 4.2e-20
C14262 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 0.0145f
C14263 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_16_7/A 0.00225f
C14264 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 3.27e-21
C14265 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 0.0215f
C14266 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_20/A 0.0137f
C14267 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_23/HI 0.00974f
C14268 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# sky130_fd_sc_hd__conb_1_47/HI 8.82e-19
C14269 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.4e-21
C14270 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.66e-20
C14271 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 1.47e-21
C14272 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__conb_1_51/HI 0.0441f
C14273 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_59/Y 0.106f
C14274 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.51e-19
C14275 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_1_29/Y 0.212f
C14276 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__conb_1_15/LO 1.71e-19
C14277 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 4.64e-19
C14278 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_647_21# -0.00122f
C14279 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# -0.00901f
C14280 V_SENSE sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 2.31e-19
C14281 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__inv_1_27/Y 2.85e-19
C14282 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# sky130_fd_sc_hd__inv_1_44/A 1.51e-19
C14283 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_3/Y 0.00964f
C14284 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 1.44e-19
C14285 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# -7.17e-20
C14286 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# -1.76e-19
C14287 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 1.78e-33
C14288 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.333f
C14289 sky130_fd_sc_hd__dfbbn_1_40/Q_N FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00229f
C14290 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_53/A 4.37e-19
C14291 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_1_19/Y 0.00149f
C14292 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__conb_1_6/HI 0.0221f
C14293 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0148f
C14294 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0168f
C14295 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0465f
C14296 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__conb_1_7/HI 0.105f
C14297 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0298f
C14298 sky130_fd_sc_hd__dfbbn_1_32/Q_N RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00881f
C14299 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__inv_1_55/Y 3.72e-19
C14300 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__conb_1_15/HI -0.00907f
C14301 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__conb_1_47/HI 7.79e-21
C14302 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.011f
C14303 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__conb_1_8/HI 0.00353f
C14304 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__conb_1_37/HI 5.77e-19
C14305 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_22/Y 3.05e-19
C14306 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1_48/Y 0.00285f
C14307 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -1.89e-19
C14308 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# -3.65e-19
C14309 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__dfbbn_1_26/Q_N 5.37e-19
C14310 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.67e-21
C14311 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 8.99e-20
C14312 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 1.07e-20
C14313 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# V_LOW 0.00556f
C14314 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# V_LOW -6.55e-19
C14315 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# V_LOW -0.0077f
C14316 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_29/LO 8.39e-19
C14317 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# V_LOW 3.56e-20
C14318 V_SENSE sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 2.31e-19
C14319 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00138f
C14320 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# V_LOW -1.01e-19
C14321 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_10/Y 2.21e-19
C14322 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00128f
C14323 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 1.01e-20
C14324 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_7/HI -0.0785f
C14325 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.28e-19
C14326 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__conb_1_9/HI 5.05e-19
C14327 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# V_LOW 0.00688f
C14328 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.27e-19
C14329 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 2.62e-21
C14330 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.0308f
C14331 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__inv_16_41/Y 0.00124f
C14332 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# V_LOW -0.00389f
C14333 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_30/HI 2.44e-19
C14334 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__conb_1_37/HI 1.08e-19
C14335 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_24/Y 5.46e-20
C14336 sky130_fd_sc_hd__inv_16_6/A RISING_COUNTER.COUNT_SUB_DFF3.Q 0.51f
C14337 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 7.06e-19
C14338 sky130_fd_sc_hd__conb_1_25/LO FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0128f
C14339 sky130_fd_sc_hd__conb_1_35/LO FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00161f
C14340 sky130_fd_sc_hd__inv_1_24/Y sky130_fd_sc_hd__inv_1_47/A 0.00388f
C14341 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__conb_1_39/HI 1.2e-19
C14342 sky130_fd_sc_hd__conb_1_14/LO FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00893f
C14343 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 0.00113f
C14344 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00869f
C14345 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# 0.00184f
C14346 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nand2_1_5/Y 4.48e-20
C14347 sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_16_2/Y 3.37e-19
C14348 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1_66/A 9.87e-21
C14349 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_1_47/Y 3.4e-21
C14350 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__dfbbn_1_0/a_27_47# 0.00388f
C14351 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_66/A 0.00277f
C14352 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 1.81e-19
C14353 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__conb_1_48/HI 5.12e-21
C14354 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__dfbbn_1_29/Q_N 1.57e-19
C14355 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 0.129f
C14356 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# V_LOW -0.00143f
C14357 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__conb_1_37/HI 0.00248f
C14358 sky130_fd_sc_hd__conb_1_41/LO V_LOW 0.0894f
C14359 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.72e-20
C14360 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# sky130_fd_sc_hd__conb_1_26/HI 4.96e-20
C14361 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# V_LOW 3.56e-20
C14362 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_55/Y 5.3e-20
C14363 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__inv_1_12/Y 0.00161f
C14364 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__inv_1_50/Y 3.33e-21
C14365 sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.75e-19
C14366 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 9.19e-19
C14367 sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__inv_1_28/Y 5.85e-22
C14368 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# sky130_fd_sc_hd__conb_1_51/HI 4.8e-19
C14369 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.22e-19
C14370 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.587f
C14371 V_SENSE sky130_fd_sc_hd__inv_16_52/A 0.347f
C14372 sky130_fd_sc_hd__conb_1_30/LO V_LOW 0.0901f
C14373 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 6.11e-20
C14374 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00243f
C14375 sky130_fd_sc_hd__inv_16_41/Y sky130_fd_sc_hd__conb_1_30/HI 0.0836f
C14376 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 0.014f
C14377 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# V_LOW -0.00266f
C14378 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# sky130_fd_sc_hd__inv_16_42/Y 2.51e-19
C14379 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.00164f
C14380 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# sky130_fd_sc_hd__conb_1_6/HI 9.26e-20
C14381 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.0429f
C14382 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_56/Y 9.9e-21
C14383 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_64/A 1.51e-20
C14384 RISING_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 1.41e-19
C14385 FULL_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0767f
C14386 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.596f
C14387 FALLING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 3.71e-20
C14388 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__conb_1_15/HI -1.41e-20
C14389 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 6.69e-19
C14390 sky130_fd_sc_hd__fill_4_215/VPB V_LOW 0.798f
C14391 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_16_19/Y 0.0719f
C14392 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_19/Y 3.02e-19
C14393 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 9.07e-19
C14394 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 1.15e-20
C14395 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# -1.76e-19
C14396 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# -5.54e-21
C14397 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -7.6e-19
C14398 sky130_fd_sc_hd__inv_1_2/Y FULL_COUNTER.COUNT_SUB_DFF6.Q 0.434f
C14399 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.72e-19
C14400 RISING_COUNTER.COUNT_SUB_DFF0.Q Reset 0.259f
C14401 sky130_fd_sc_hd__nand2_8_4/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00566f
C14402 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/Q_N 2.1e-19
C14403 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# 6.96e-19
C14404 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_46/A 0.256f
C14405 sky130_fd_sc_hd__inv_16_23/A sky130_fd_sc_hd__inv_16_20/A 0.0906f
C14406 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_64/A 0.0771f
C14407 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_473_413# -0.0103f
C14408 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# -0.00224f
C14409 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 6.31e-21
C14410 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# 3.23e-21
C14411 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF8.Q 5.8e-19
C14412 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0373f
C14413 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__conb_1_37/HI 1.69e-19
C14414 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__nor2_1_0/Y 1.38e-21
C14415 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__conb_1_0/HI 1.31e-19
C14416 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_1_23/A 6.61e-19
C14417 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 0.0226f
C14418 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# sky130_fd_sc_hd__conb_1_39/HI 1.27e-20
C14419 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00217f
C14420 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_58/Y 0.0296f
C14421 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 0.00275f
C14422 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__conb_1_24/HI 3.09e-19
C14423 sky130_fd_sc_hd__conb_1_20/LO sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 0.00169f
C14424 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00511f
C14425 sky130_fd_sc_hd__conb_1_43/LO V_LOW 0.0808f
C14426 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__inv_1_13/Y 1.49e-19
C14427 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0223f
C14428 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_50/HI 0.00897f
C14429 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 9.46e-20
C14430 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# -0.00263f
C14431 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -7.6e-19
C14432 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# -5.54e-21
C14433 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0822f
C14434 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 0.00291f
C14435 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 1.73e-19
C14436 FALLING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 1.58e-21
C14437 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_53/Y 0.00595f
C14438 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 5.36e-19
C14439 sky130_fd_sc_hd__conb_1_32/LO V_LOW 0.094f
C14440 sky130_fd_sc_hd__inv_16_26/Y sky130_fd_sc_hd__inv_16_7/A 7.73e-19
C14441 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_1_22/Y 4.81e-21
C14442 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.8e-19
C14443 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 3.13e-21
C14444 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 7.72e-21
C14445 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.62e-19
C14446 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 7.41e-19
C14447 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__conb_1_44/HI 2.43e-19
C14448 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__conb_1_48/HI 1.36e-19
C14449 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_26/HI 0.314f
C14450 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# V_LOW -0.00121f
C14451 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q -1.27e-20
C14452 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 3e-20
C14453 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00454f
C14454 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00451f
C14455 sky130_fd_sc_hd__inv_16_29/A V_LOW 0.224f
C14456 sky130_fd_sc_hd__inv_1_59/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 3.17e-21
C14457 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__inv_16_42/Y 0.0119f
C14458 sky130_fd_sc_hd__dfbbn_1_42/a_581_47# sky130_fd_sc_hd__inv_16_42/Y 0.00179f
C14459 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__conb_1_37/HI 1.26e-19
C14460 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_16_41/Y 0.0294f
C14461 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_16_42/Y 0.117f
C14462 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_26/HI 0.0259f
C14463 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__conb_1_27/HI 0.322f
C14464 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00141f
C14465 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 1.99e-19
C14466 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 1.19e-19
C14467 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 1.19e-19
C14468 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 1.99e-19
C14469 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 2.11e-19
C14470 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 6.38e-19
C14471 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.0228f
C14472 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 2.11e-19
C14473 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 6.38e-19
C14474 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_31/HI 1.07e-19
C14475 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_647_21# -0.00499f
C14476 sky130_fd_sc_hd__inv_16_26/A V_LOW 0.242f
C14477 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.00159f
C14478 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_1_0/Y 0.0446f
C14479 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__inv_16_42/Y 0.0398f
C14480 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# V_LOW -0.00412f
C14481 sky130_fd_sc_hd__inv_1_37/Y sky130_fd_sc_hd__conb_1_32/LO 5.94e-19
C14482 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.91e-19
C14483 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__conb_1_15/HI -2.17e-19
C14484 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 3.4e-20
C14485 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# -2.37e-19
C14486 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# -3.07e-19
C14487 sky130_fd_sc_hd__inv_16_5/A sky130_fd_sc_hd__inv_16_7/A 0.0245f
C14488 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 9.65e-21
C14489 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__conb_1_46/HI 0.446f
C14490 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_24/A 6.59e-19
C14491 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__conb_1_35/HI 0.0431f
C14492 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.58e-19
C14493 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 1.54e-20
C14494 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.88e-20
C14495 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__conb_1_40/HI -1.6e-19
C14496 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 5.44e-20
C14497 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 4.48e-19
C14498 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_68/Y 0.00298f
C14499 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__conb_1_46/HI 8.68e-20
C14500 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_40/Y 0.308f
C14501 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# V_LOW 1.38e-19
C14502 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 1.13e-19
C14503 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 9.54e-19
C14504 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 0.00108f
C14505 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 4.99e-19
C14506 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# -0.00125f
C14507 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_381_47# -4.5e-20
C14508 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# -9.41e-19
C14509 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_16_19/Y 2.02e-19
C14510 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 7.66e-20
C14511 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand2_1_5/Y 5.91e-21
C14512 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.00996f
C14513 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 3.58e-19
C14514 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_45/Y 0.00135f
C14515 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.206f
C14516 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__inv_1_7/Y 0.00627f
C14517 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0.0269f
C14518 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 8.44e-19
C14519 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00146f
C14520 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__conb_1_37/HI 0.0075f
C14521 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 0.00104f
C14522 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 0.00215f
C14523 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 0.0112f
C14524 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__inv_1_26/Y 5.98e-19
C14525 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 1.17e-19
C14526 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__inv_16_40/Y 0.00726f
C14527 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# FULL_COUNTER.COUNT_SUB_DFF12.Q 7e-19
C14528 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# sky130_fd_sc_hd__conb_1_24/HI 0.00183f
C14529 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.52e-19
C14530 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_16_41/Y 0.561f
C14531 sky130_fd_sc_hd__inv_1_68/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00502f
C14532 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 4.8e-19
C14533 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.00318f
C14534 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_27/HI 2.86e-19
C14535 sky130_fd_sc_hd__conb_1_26/HI sky130_fd_sc_hd__inv_1_31/Y 0.294f
C14536 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_64/A 0.102f
C14537 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# V_LOW 0.0159f
C14538 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0217f
C14539 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__nand2_1_2/A 5.7e-19
C14540 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__conb_1_9/HI -6.68e-21
C14541 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# -9.32e-20
C14542 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# -4.66e-20
C14543 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# -3.79e-20
C14544 sky130_fd_sc_hd__conb_1_45/HI V_LOW 0.0313f
C14545 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 1.34e-19
C14546 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.01f
C14547 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.22e-20
C14548 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_16_40/Y 1.92e-20
C14549 sky130_fd_sc_hd__nand3_1_1/a_193_47# sky130_fd_sc_hd__inv_1_66/Y 0.00133f
C14550 sky130_fd_sc_hd__conb_1_3/LO FULL_COUNTER.COUNT_SUB_DFF6.Q 0.0109f
C14551 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.8e-20
C14552 sky130_fd_sc_hd__fill_8_949/VPB V_LOW 0.797f
C14553 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# sky130_fd_sc_hd__inv_1_39/Y 6.86e-20
C14554 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0174f
C14555 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__inv_1_22/Y 1.38e-20
C14556 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.14e-19
C14557 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.96e-20
C14558 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__conb_1_14/HI 0.0124f
C14559 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__conb_1_48/HI -6.57e-19
C14560 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0177f
C14561 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 1.01e-21
C14562 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 1.11e-20
C14563 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_47/A 1.93e-20
C14564 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 6.15e-20
C14565 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_39/HI -0.0499f
C14566 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__inv_16_42/Y 0.00576f
C14567 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 3.87e-19
C14568 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1_44/HI 0.0457f
C14569 sky130_fd_sc_hd__inv_16_3/A sky130_fd_sc_hd__inv_16_28/Y 0.00176f
C14570 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__inv_1_50/Y 0.00131f
C14571 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# sky130_fd_sc_hd__inv_16_42/Y 6.53e-19
C14572 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_1_31/Y 3.03e-19
C14573 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_8/A 0.064f
C14574 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_30/Y 0.62f
C14575 Reset FULL_COUNTER.COUNT_SUB_DFF1.Q 1.37f
C14576 sky130_fd_sc_hd__nand2_8_4/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0198f
C14577 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_48/a_791_47# -0.0121f
C14578 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 0.0126f
C14579 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_581_47# -2.6e-20
C14580 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00983f
C14581 sky130_fd_sc_hd__conb_1_29/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.201f
C14582 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_16_40/Y 8.07e-20
C14583 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# sky130_fd_sc_hd__inv_16_42/Y 0.00482f
C14584 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# V_LOW -1.39e-35
C14585 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# -1.66e-19
C14586 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# -7.17e-20
C14587 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_25/LO 4.48e-21
C14588 sky130_fd_sc_hd__inv_1_48/Y V_LOW 0.0917f
C14589 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__inv_1_59/Y 0.0386f
C14590 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/Q_N -4.33e-20
C14591 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__nand3_1_2/Y 2.04e-20
C14592 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# sky130_fd_sc_hd__conb_1_35/HI 4.99e-19
C14593 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 7.09e-21
C14594 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# sky130_fd_sc_hd__conb_1_40/HI -0.00125f
C14595 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0061f
C14596 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00126f
C14597 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.0323f
C14598 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__conb_1_46/HI 1.04e-19
C14599 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__inv_16_40/Y 0.0471f
C14600 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.98e-19
C14601 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# V_LOW 4.8e-20
C14602 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# -1.69e-19
C14603 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# -0.0103f
C14604 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -5.84e-19
C14605 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_1_49/Y 3.73e-20
C14606 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# 1.16e-19
C14607 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 4.57e-21
C14608 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00134f
C14609 sky130_fd_sc_hd__conb_1_0/LO FULL_COUNTER.COUNT_SUB_DFF6.Q 2.96e-19
C14610 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 4.49e-21
C14611 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 7.44e-21
C14612 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 4.58e-19
C14613 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 2.38e-20
C14614 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# 0.00146f
C14615 V_SENSE sky130_fd_sc_hd__conb_1_47/LO 9.19e-19
C14616 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_19/A 0.00223f
C14617 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 5.69e-20
C14618 V_SENSE FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0946f
C14619 FALLING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.23e-19
C14620 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__conb_1_51/HI 2.68e-19
C14621 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__inv_1_32/Y 3.43e-21
C14622 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 3.99e-19
C14623 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 0.0104f
C14624 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.74e-20
C14625 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 5.23e-20
C14626 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_16_41/Y 0.0672f
C14627 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__inv_16_40/Y 0.0313f
C14628 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# sky130_fd_sc_hd__inv_1_2/Y 5.11e-19
C14629 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# V_LOW 1.38e-19
C14630 sky130_fd_sc_hd__inv_16_40/Y FULL_COUNTER.COUNT_SUB_DFF0.Q 0.29f
C14631 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_30/HI 2.53e-20
C14632 sky130_fd_sc_hd__inv_1_18/A sky130_fd_sc_hd__inv_16_2/Y 6.69e-20
C14633 sky130_fd_sc_hd__inv_1_66/A V_LOW 0.34f
C14634 sky130_fd_sc_hd__inv_1_58/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 0.125f
C14635 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# 1.07e-21
C14636 sky130_fd_sc_hd__inv_16_48/Y sky130_fd_sc_hd__inv_16_51/Y 2.46f
C14637 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_891_329# -2.2e-20
C14638 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# -0.00161f
C14639 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0334f
C14640 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# V_LOW 0.00478f
C14641 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00115f
C14642 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# sky130_fd_sc_hd__conb_1_9/HI 1.24e-20
C14643 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.45e-20
C14644 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/Q_N -4.33e-20
C14645 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__conb_1_3/HI -0.00907f
C14646 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_1_34/Y 3.76e-21
C14647 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# V_LOW 0.0145f
C14648 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_44/A 7.36e-20
C14649 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00337f
C14650 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.154f
C14651 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00354f
C14652 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.61e-19
C14653 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__inv_16_41/Y 0.0824f
C14654 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_1_11/Y 6.27e-19
C14655 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# sky130_fd_sc_hd__conb_1_14/HI -0.00257f
C14656 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_9/Y 1.66e-19
C14657 sky130_fd_sc_hd__conb_1_27/HI V_LOW 0.373f
C14658 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.022f
C14659 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__nand3_1_2/Y 4.29e-19
C14660 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# 0.0141f
C14661 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 7.81e-20
C14662 sky130_fd_sc_hd__inv_1_0/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 7.39e-19
C14663 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.311f
C14664 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00162f
C14665 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_8/LO 3.08e-20
C14666 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_27/Y 0.0257f
C14667 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.85e-21
C14668 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# Reset 6.92e-19
C14669 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_23/HI 0.0228f
C14670 RISING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF14.Q 2.14f
C14671 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 7.85e-21
C14672 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0.00219f
C14673 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 1.82e-20
C14674 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 3.05e-22
C14675 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 2.6e-20
C14676 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.74e-20
C14677 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__inv_16_41/Y 2.97e-20
C14678 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0161f
C14679 sky130_fd_sc_hd__dfbbn_1_23/Q_N V_LOW -0.00993f
C14680 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# sky130_fd_sc_hd__conb_1_2/HI 2.05e-19
C14681 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00261f
C14682 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# -0.134f
C14683 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__conb_1_26/HI 3.65e-20
C14684 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_25/HI 1.02e-20
C14685 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0145f
C14686 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.82e-20
C14687 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_28/Y 0.072f
C14688 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_1_21/Y 0.0296f
C14689 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# 2.75e-19
C14690 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_581_47# -7.91e-19
C14691 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__inv_1_1/Y 7.85e-22
C14692 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# -6.8e-19
C14693 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 7.71e-21
C14694 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 1.48e-20
C14695 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__inv_1_49/Y 6.08e-21
C14696 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.84e-19
C14697 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__conb_1_10/HI 0.027f
C14698 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/Q_N 7.69e-19
C14699 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/Q_N -9.56e-20
C14700 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_1_40/Y 1.19e-20
C14701 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.86e-19
C14702 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.29e-20
C14703 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# -4.66e-20
C14704 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# -3.79e-20
C14705 sky130_fd_sc_hd__conb_1_9/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.123f
C14706 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# sky130_fd_sc_hd__inv_1_3/Y 3.75e-21
C14707 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__dfbbn_1_40/a_473_413# 6.86e-21
C14708 sky130_fd_sc_hd__inv_16_52/A CLOCK_GEN.SR_Op.Q 0.034f
C14709 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__conb_1_51/HI 2.38e-19
C14710 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 1.95e-20
C14711 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 9.98e-20
C14712 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 5.34e-19
C14713 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 6.48e-20
C14714 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 6.63e-20
C14715 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 3.1e-20
C14716 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_16_41/Y 0.0528f
C14717 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 1.24e-19
C14718 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 4.12e-20
C14719 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# -0.00149f
C14720 FULL_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0331f
C14721 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__inv_16_41/Y 0.00432f
C14722 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# V_LOW -0.01f
C14723 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# V_LOW -0.312f
C14724 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# V_LOW 3.56e-20
C14725 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# -3.46e-20
C14726 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_557_413# -3.67e-20
C14727 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# -6.29e-19
C14728 sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__conb_1_9/HI 4.59e-21
C14729 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 5.61e-19
C14730 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# sky130_fd_sc_hd__conb_1_3/HI -9.71e-19
C14731 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/Q_N -2.84e-32
C14732 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# sky130_fd_sc_hd__inv_1_60/Y 2.63e-19
C14733 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_31/Y 0.167f
C14734 sky130_fd_sc_hd__inv_1_44/A FULL_COUNTER.COUNT_SUB_DFF1.Q 0.179f
C14735 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.686f
C14736 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_891_329# -2.2e-20
C14737 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# -3.48e-20
C14738 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# sky130_fd_sc_hd__inv_16_41/Y 5.14e-21
C14739 sky130_fd_sc_hd__inv_1_61/Y V_LOW 0.0155f
C14740 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# sky130_fd_sc_hd__inv_16_40/Y 0.00644f
C14741 FULL_COUNTER.COUNT_SUB_DFF16.Q V_LOW 2.96f
C14742 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0356f
C14743 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# 5.57e-19
C14744 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 6.94e-19
C14745 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 0.0331f
C14746 sky130_fd_sc_hd__inv_1_1/Y V_LOW 0.19f
C14747 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__inv_1_29/Y 3.86e-19
C14748 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__conb_1_26/HI 0.0341f
C14749 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 0.00782f
C14750 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# 2.59e-19
C14751 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 0.00116f
C14752 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0.00126f
C14753 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_12/Q_N 6.01e-21
C14754 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_16_40/Y 0.0342f
C14755 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 3.29e-20
C14756 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__inv_1_9/Y 5.21e-21
C14757 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__conb_1_8/LO 5.6e-20
C14758 sky130_fd_sc_hd__nor2_1_0/a_109_297# V_LOW -0.002f
C14759 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__conb_1_31/HI 1.5e-19
C14760 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 1.96e-20
C14761 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.96e-21
C14762 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 2.81e-21
C14763 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 1.96e-20
C14764 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 4.58e-19
C14765 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nand2_8_9/A 0.00164f
C14766 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 3.14e-19
C14767 sky130_fd_sc_hd__inv_16_24/Y sky130_fd_sc_hd__inv_16_22/A 0.00855f
C14768 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# -3.79e-20
C14769 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# -4.66e-20
C14770 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_1_32/Y 0.00211f
C14771 sky130_fd_sc_hd__conb_1_25/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0329f
C14772 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# V_LOW 0.015f
C14773 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_28/Y 0.0309f
C14774 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 1.07e-20
C14775 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 2.29e-19
C14776 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 0.0134f
C14777 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# sky130_fd_sc_hd__inv_1_69/Y 4.29e-21
C14778 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.00245f
C14779 sky130_fd_sc_hd__inv_1_59/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0261f
C14780 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 7.35e-19
C14781 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00182f
C14782 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 5.79e-19
C14783 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__dfbbn_1_43/a_891_329# 0.00127f
C14784 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_1_36/Y 9.72e-22
C14785 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00291f
C14786 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__inv_1_50/Y 6.64e-20
C14787 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0.0211f
C14788 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# -0.0571f
C14789 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.6e-20
C14790 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 3.33e-19
C14791 sky130_fd_sc_hd__dfbbn_1_28/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 1.89e-19
C14792 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__inv_16_41/Y 0.0633f
C14793 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 0.0196f
C14794 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# V_LOW 0.0121f
C14795 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_1_36/Y 2.25e-21
C14796 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_16_40/Y 0.0129f
C14797 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# 1.05e-19
C14798 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_581_47# -2.6e-20
C14799 sky130_fd_sc_hd__conb_1_34/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 9.11e-19
C14800 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_47/Y 3.01e-19
C14801 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__inv_16_41/Y 0.00558f
C14802 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# V_LOW -6.55e-19
C14803 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__inv_1_33/Y 0.0315f
C14804 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_1_35/Y 3.5e-20
C14805 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 1.28e-19
C14806 sky130_fd_sc_hd__inv_8_0/A sky130_fd_sc_hd__inv_16_2/Y 0.0487f
C14807 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# V_LOW 4.8e-20
C14808 sky130_fd_sc_hd__dfbbn_1_48/Q_N FALLING_COUNTER.COUNT_SUB_DFF4.Q 3.21e-19
C14809 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -7.6e-19
C14810 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# -5.54e-21
C14811 sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__conb_1_3/HI -2.17e-19
C14812 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# Reset 0.00142f
C14813 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# sky130_fd_sc_hd__inv_1_44/A 2.24e-19
C14814 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# -0.00196f
C14815 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# V_LOW 2.26e-20
C14816 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.128f
C14817 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.35e-19
C14818 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# V_LOW 0.0137f
C14819 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 6.09e-21
C14820 sky130_fd_sc_hd__conb_1_39/HI CLOCK_GEN.SR_Op.Q 2.74e-19
C14821 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.04f
C14822 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_25/HI 1.85e-20
C14823 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__nor2_1_0/Y 4.43e-20
C14824 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__conb_1_37/HI 2.15e-20
C14825 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00345f
C14826 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__inv_16_40/Y 2.48e-20
C14827 FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00365f
C14828 V_SENSE sky130_fd_sc_hd__inv_16_27/Y 0.146f
C14829 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_193_47# -0.206f
C14830 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 1.25e-19
C14831 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 1.25e-19
C14832 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 7.69e-20
C14833 FALLING_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0289f
C14834 sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__inv_1_66/A 5.55e-19
C14835 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.00106f
C14836 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.0029f
C14837 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.0035f
C14838 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__conb_1_35/LO 0.00434f
C14839 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.3e-19
C14840 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__conb_1_34/HI 5.9e-22
C14841 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/Q_N 6.91e-19
C14842 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 1.12e-20
C14843 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 1.44e-20
C14844 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__inv_1_43/Y 0.00211f
C14845 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00299f
C14846 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_12/LO 4.33e-21
C14847 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__nand2_1_1/a_113_47# 1.84e-20
C14848 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__inv_16_40/Y 0.0391f
C14849 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_24/Y 1.79e-19
C14850 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 0.0107f
C14851 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00225f
C14852 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__nand2_1_5/Y 4.22e-19
C14853 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# -6.43e-20
C14854 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# -3.06e-20
C14855 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__conb_1_31/HI 1.92e-20
C14856 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# V_LOW 4.8e-20
C14857 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.74e-19
C14858 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_1_8/Y 0.00702f
C14859 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.00172f
C14860 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__inv_1_12/Y 6.45e-20
C14861 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 6.42e-21
C14862 sky130_fd_sc_hd__conb_1_32/HI RISING_COUNTER.COUNT_SUB_DFF8.Q 0.101f
C14863 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# V_LOW 0.0258f
C14864 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 3.08e-20
C14865 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 3.61e-20
C14866 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 2.09e-19
C14867 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_26/HI 0.0212f
C14868 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00263f
C14869 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 0.194f
C14870 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# V_LOW 1.79e-20
C14871 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__inv_1_28/Y 0.00574f
C14872 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 9.69e-21
C14873 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_64/A 0.00246f
C14874 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF14.Q 4.18e-19
C14875 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 8.6e-20
C14876 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# 1.86e-21
C14877 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# 9.18e-21
C14878 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# V_LOW 0.0156f
C14879 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF2.Q 0.0169f
C14880 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 4.57e-19
C14881 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__inv_1_24/Y 7.17e-21
C14882 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_16_42/Y 0.366f
C14883 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__conb_1_47/HI 0.00541f
C14884 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_47/A 5.69e-19
C14885 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# 3.5e-19
C14886 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# 7.51e-21
C14887 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00493f
C14888 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# -1.24e-20
C14889 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.82e-20
C14890 sky130_fd_sc_hd__conb_1_0/HI FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0234f
C14891 Reset FULL_COUNTER.COUNT_SUB_DFF0.Q 2.74f
C14892 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# sky130_fd_sc_hd__inv_16_41/Y 0.00501f
C14893 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF2.Q 6.06e-19
C14894 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# V_LOW -0.00728f
C14895 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__inv_16_40/Y 7.23e-20
C14896 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_1_35/Y 2.64e-20
C14897 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__inv_16_41/Y 0.00463f
C14898 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0024f
C14899 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_16_40/Y 6.97e-22
C14900 V_SENSE sky130_fd_sc_hd__inv_1_52/A 2.01e-19
C14901 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# V_LOW -0.107f
C14902 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF14.Q 1.44e-19
C14903 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF15.Q 7.13e-22
C14904 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_16_2/Y 0.178f
C14905 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# -4.1e-19
C14906 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_891_329# -2.2e-20
C14907 sky130_fd_sc_hd__nand2_1_0/a_113_47# V_LOW -1.78e-19
C14908 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_8/HI 0.0244f
C14909 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 3.24e-22
C14910 sky130_fd_sc_hd__conb_1_45/LO FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.003f
C14911 sky130_fd_sc_hd__inv_16_42/Y sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 2.76e-20
C14912 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.38e-20
C14913 sky130_fd_sc_hd__dfbbn_1_25/Q_N FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0233f
C14914 V_SENSE sky130_fd_sc_hd__inv_16_51/Y 6.95f
C14915 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 0.00106f
C14916 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_19/Q_N 0.026f
C14917 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_34/HI 0.00137f
C14918 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 5.74e-20
C14919 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__conb_1_34/HI 8.31e-20
C14920 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 9.3e-22
C14921 sky130_fd_sc_hd__inv_16_23/Y sky130_fd_sc_hd__inv_16_20/A 0.0309f
C14922 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_32/Y 0.222f
C14923 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/Q_N 9.64e-20
C14924 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 0.028f
C14925 FULL_COUNTER.COUNT_SUB_DFF2.Q CLOCK_GEN.SR_Op.Q 0.0221f
C14926 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF8.Q 1.02e-20
C14927 sky130_fd_sc_hd__inv_16_50/Y sky130_fd_sc_hd__inv_16_50/A 0.0399f
C14928 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# sky130_fd_sc_hd__conb_1_30/HI 0.00138f
C14929 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_2_0/A 3.35e-20
C14930 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_41/Y 5.98e-20
C14931 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_19/HI -0.00398f
C14932 sky130_fd_sc_hd__inv_16_6/A sky130_fd_sc_hd__conb_1_35/HI 0.00112f
C14933 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 3.7e-19
C14934 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 2.01e-19
C14935 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 2.01e-19
C14936 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 3.7e-19
C14937 sky130_fd_sc_hd__inv_1_58/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.173f
C14938 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.028f
C14939 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 0.00319f
C14940 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__conb_1_28/LO 0.0015f
C14941 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__conb_1_21/HI 0.0116f
C14942 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# V_LOW 2.94e-20
C14943 sky130_fd_sc_hd__nand2_8_2/a_27_47# V_LOW -0.00644f
C14944 sky130_fd_sc_hd__conb_1_31/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.503f
C14945 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0.00184f
C14946 sky130_fd_sc_hd__inv_16_47/Y sky130_fd_sc_hd__inv_16_51/A 5.81f
C14947 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_1_64/A 1.56e-19
C14948 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF12.Q 3.18e-19
C14949 sky130_fd_sc_hd__dfbbn_1_50/a_581_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.86e-19
C14950 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 2.04e-20
C14951 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.73e-20
C14952 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# V_LOW -3.52e-20
C14953 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_22/Y 0.00129f
C14954 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__inv_1_62/Y 0.086f
C14955 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_891_329# -0.00159f
C14956 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# -0.00851f
C14957 sky130_fd_sc_hd__conb_1_47/LO sky130_fd_sc_hd__inv_1_63/Y 0.00179f
C14958 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# V_LOW -9.15e-19
C14959 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00597f
C14960 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 8.66e-21
C14961 FULL_COUNTER.COUNT_SUB_DFF17.Q V_LOW 1.47f
C14962 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF8.Q 0.00286f
C14963 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__inv_1_50/Y 1.17e-19
C14964 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_581_47# -2.6e-20
C14965 FALLING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 0.533f
C14966 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_66/Y 0.263f
C14967 sky130_fd_sc_hd__inv_16_42/Y V_LOW 1.58f
C14968 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__inv_1_35/Y 2.66e-21
C14969 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_16_40/Y 0.00355f
C14970 V_SENSE sky130_fd_sc_hd__inv_1_46/A 0.615f
C14971 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__nand3_1_2/Y 1.63e-19
C14972 sky130_fd_sc_hd__inv_1_24/Y Reset 0.0554f
C14973 sky130_fd_sc_hd__conb_1_49/LO V_LOW 0.138f
C14974 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# V_LOW 0.006f
C14975 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__inv_16_40/Y 2.33e-19
C14976 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# -0.00631f
C14977 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# -0.00988f
C14978 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# V_LOW -2.68e-19
C14979 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# -0.00385f
C14980 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/Q_N -4.78e-20
C14981 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# sky130_fd_sc_hd__inv_1_41/Y 5.11e-19
C14982 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__conb_1_8/HI 0.00616f
C14983 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 4.69e-21
C14984 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__conb_1_35/HI 7.72e-22
C14985 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# -0.00631f
C14986 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# -0.00591f
C14987 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 1.25e-20
C14988 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI 8.83e-19
C14989 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_66/A 2.8e-19
C14990 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__conb_1_35/HI 6.59e-20
C14991 sky130_fd_sc_hd__inv_1_56/Y sky130_fd_sc_hd__inv_1_64/A 4.69e-20
C14992 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__conb_1_17/HI 0.0131f
C14993 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00364f
C14994 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_27/HI -0.00154f
C14995 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# sky130_fd_sc_hd__conb_1_34/HI -0.00246f
C14996 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__conb_1_38/HI 1.62e-19
C14997 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_25/Y -0.00409f
C14998 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_16_42/Y 2.27e-20
C14999 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__conb_1_20/HI 0.00535f
C15000 sky130_fd_sc_hd__conb_1_9/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.17f
C15001 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 2.42e-19
C15002 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_26/Y 1.21e-19
C15003 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# 3.94e-20
C15004 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_381_47# -0.00833f
C15005 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# -0.00117f
C15006 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__conb_1_19/HI 0.00126f
C15007 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0018f
C15008 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0386f
C15009 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# -2.52e-19
C15010 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# -0.00151f
C15011 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0192f
C15012 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_25/LO 8.84e-20
C15013 sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__inv_16_41/Y 0.601f
C15014 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0151f
C15015 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__inv_1_34/Y 0.0141f
C15016 RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 2.11e-20
C15017 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 2.96f
C15018 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 1.79e-20
C15019 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 1.79e-20
C15020 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_69/Y 0.588f
C15021 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 2.04e-19
C15022 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 6.62e-21
C15023 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 9.12e-19
C15024 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.00124f
C15025 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00635f
C15026 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_29/Y 6.96e-20
C15027 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.0126f
C15028 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 6.81e-19
C15029 sky130_fd_sc_hd__inv_1_44/A FULL_COUNTER.COUNT_SUB_DFF0.Q 0.0286f
C15030 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__inv_1_31/Y 1.82e-20
C15031 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_10/HI 2.17e-20
C15032 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0.00315f
C15033 sky130_fd_sc_hd__inv_1_65/A sky130_fd_sc_hd__inv_1_67/A 7.15e-21
C15034 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__inv_1_38/Y 2.72e-19
C15035 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.22e-19
C15036 V_LOW V_GND 2.3p
C15037 FULL_COUNTER.COUNT_SUB_DFF16.Q V_GND 4.18f
C15038 FULL_COUNTER.COUNT_SUB_DFF14.Q V_GND 5.68f
C15039 FULL_COUNTER.COUNT_SUB_DFF13.Q V_GND 4.89f
C15040 RISING_COUNTER.COUNT_SUB_DFF10.Q V_GND 1.87f
C15041 FALLING_COUNTER.COUNT_SUB_DFF9.Q V_GND 1.32f
C15042 RISING_COUNTER.COUNT_SUB_DFF8.Q V_GND 4.43f
C15043 FULL_COUNTER.COUNT_SUB_DFF12.Q V_GND 5.03f
C15044 FULL_COUNTER.COUNT_SUB_DFF11.Q V_GND 4.03f
C15045 FULL_COUNTER.COUNT_SUB_DFF10.Q V_GND 2.89f
C15046 RISING_COUNTER.COUNT_SUB_DFF6.Q V_GND 3.3f
C15047 FALLING_COUNTER.COUNT_SUB_DFF5.Q V_GND 3.89f
C15048 RISING_COUNTER.COUNT_SUB_DFF5.Q V_GND 7.39f
C15049 FULL_COUNTER.COUNT_SUB_DFF9.Q V_GND 3.78f
C15050 RISING_COUNTER.COUNT_SUB_DFF4.Q V_GND 4.49f
C15051 FALLING_COUNTER.COUNT_SUB_DFF3.Q V_GND 3.25f
C15052 FULL_COUNTER.COUNT_SUB_DFF8.Q V_GND 3.92f
C15053 RISING_COUNTER.COUNT_SUB_DFF3.Q V_GND 6.91f
C15054 FULL_COUNTER.COUNT_SUB_DFF7.Q V_GND 3.85f
C15055 FULL_COUNTER.COUNT_SUB_DFF5.Q V_GND 2.93f
C15056 FALLING_COUNTER.COUNT_SUB_DFF0.Q V_GND 7.27f
C15057 FULL_COUNTER.COUNT_SUB_DFF1.Q V_GND 4.91f
C15058 FULL_COUNTER.COUNT_SUB_DFF0.Q V_GND 6.95f
C15059 CLOCK_GEN.SR_Op.Q V_GND 4.91f
C15060 V_HIGH V_GND 0.614p
C15061 FULL_COUNTER.COUNT_SUB_DFF17.Q V_GND 5.76f
C15062 sky130_fd_sc_hd__conb_1_11/HI V_GND 0.5f
C15063 FULL_COUNTER.COUNT_SUB_DFF18.Q V_GND 8.31f
C15064 sky130_fd_sc_hd__conb_1_15/HI V_GND 0.638f
C15065 sky130_fd_sc_hd__conb_1_16/HI V_GND 0.319f
C15066 sky130_fd_sc_hd__inv_1_27/Y V_GND 0.349f
C15067 sky130_fd_sc_hd__conb_1_19/HI V_GND 0.656f
C15068 sky130_fd_sc_hd__conb_1_17/HI V_GND 0.69f
C15069 sky130_fd_sc_hd__inv_1_26/Y V_GND 0.352f
C15070 sky130_fd_sc_hd__conb_1_23/HI V_GND 0.378f
C15071 sky130_fd_sc_hd__inv_1_31/Y V_GND 0.199f
C15072 sky130_fd_sc_hd__conb_1_26/HI V_GND 0.983f
C15073 sky130_fd_sc_hd__inv_1_29/Y V_GND 0.632f
C15074 sky130_fd_sc_hd__inv_1_28/Y V_GND 0.334f
C15075 sky130_fd_sc_hd__inv_1_30/Y V_GND 0.303f
C15076 sky130_fd_sc_hd__inv_1_58/Y V_GND 0.484f
C15077 sky130_fd_sc_hd__conb_1_30/HI V_GND 0.611f
C15078 sky130_fd_sc_hd__inv_1_38/Y V_GND 0.32f
C15079 sky130_fd_sc_hd__inv_1_40/Y V_GND 0.192f
C15080 sky130_fd_sc_hd__conb_1_8/HI V_GND 0.374f
C15081 sky130_fd_sc_hd__inv_16_41/Y V_GND 14.6f
C15082 sky130_fd_sc_hd__conb_1_32/HI V_GND 0.593f
C15083 sky130_fd_sc_hd__inv_1_10/Y V_GND 1f
C15084 sky130_fd_sc_hd__conb_1_6/HI V_GND 0.545f
C15085 sky130_fd_sc_hd__inv_1_35/Y V_GND 0.151f
C15086 sky130_fd_sc_hd__conb_1_29/HI V_GND 0.748f
C15087 sky130_fd_sc_hd__inv_1_41/Y V_GND 0.323f
C15088 sky130_fd_sc_hd__conb_1_27/HI V_GND 0.422f
C15089 sky130_fd_sc_hd__inv_1_59/Y V_GND 0.34f
C15090 FALLING_COUNTER.COUNT_SUB_DFF6.Q V_GND 3.84f
C15091 FALLING_COUNTER.COUNT_SUB_DFF4.Q V_GND 5.28f
C15092 sky130_fd_sc_hd__inv_1_39/Y V_GND 0.303f
C15093 sky130_fd_sc_hd__conb_1_38/HI V_GND 0.644f
C15094 sky130_fd_sc_hd__inv_1_49/Y V_GND 0.322f
C15095 sky130_fd_sc_hd__conb_1_40/HI V_GND 0.473f
C15096 sky130_fd_sc_hd__conb_1_2/HI V_GND 0.483f
C15097 sky130_fd_sc_hd__inv_1_1/Y V_GND 0.216f
C15098 sky130_fd_sc_hd__inv_1_45/Y V_GND 0.449f
C15099 sky130_fd_sc_hd__inv_1_48/Y V_GND 0.977f
C15100 sky130_fd_sc_hd__conb_1_37/HI V_GND 0.386f
C15101 sky130_fd_sc_hd__inv_1_64/Y V_GND 0.355f
C15102 sky130_fd_sc_hd__inv_1_64/A V_GND 0.989f
C15103 sky130_fd_sc_hd__inv_1_56/Y V_GND 0.697f
C15104 sky130_fd_sc_hd__inv_1_44/A V_GND 0.818f
C15105 transmission_gate_9/GN V_GND 4.73f
C15106 Reset V_GND 36.1f
C15107 sky130_fd_sc_hd__inv_16_2/Y V_GND 4.74f
C15108 sky130_fd_sc_hd__inv_1_47/Y V_GND 0.703f
C15109 sky130_fd_sc_hd__inv_1_66/A V_GND 2.29f
C15110 sky130_fd_sc_hd__nand2_1_5/Y V_GND 0.182f
C15111 sky130_fd_sc_hd__inv_1_19/Y V_GND 0.9f
C15112 sky130_fd_sc_hd__inv_16_8/Y V_GND 1.45f
C15113 sky130_fd_sc_hd__inv_16_8/A V_GND 1.49f
C15114 sky130_fd_sc_hd__inv_16_9/Y V_GND 1.57f
C15115 sky130_fd_sc_hd__inv_16_28/Y V_GND 1.53f
C15116 sky130_fd_sc_hd__inv_1_67/A V_GND 2.56f
C15117 sky130_fd_sc_hd__inv_16_29/A V_GND 1.47f
C15118 sky130_fd_sc_hd__inv_1_24/A V_GND 1.97f
C15119 sky130_fd_sc_hd__inv_16_22/A V_GND 1.73f
C15120 sky130_fd_sc_hd__inv_16_29/Y V_GND 1.69f
C15121 sky130_fd_sc_hd__inv_16_24/Y V_GND 1.85f
C15122 sky130_fd_sc_hd__inv_16_32/Y V_GND 1.72f
C15123 sky130_fd_sc_hd__inv_16_15/A V_GND 1.72f
C15124 sky130_fd_sc_hd__inv_16_15/Y V_GND 1.51f
C15125 sky130_fd_sc_hd__inv_16_50/A V_GND 3.42f
C15126 sky130_fd_sc_hd__inv_16_48/A V_GND 5.82f
C15127 sky130_fd_sc_hd__inv_16_55/Y V_GND 1.59f
C15128 sky130_fd_sc_hd__inv_16_51/Y V_GND 1.93f
C15129 sky130_fd_sc_hd__inv_16_49/A V_GND 8.4f
C15130 sky130_fd_sc_hd__inv_16_51/A V_GND 6.22f
C15131 sky130_fd_sc_hd__inv_16_47/Y V_GND 6.54f
C15132 FULL_COUNTER.COUNT_SUB_DFF6.Q V_GND 3.4f
C15133 sky130_fd_sc_hd__inv_1_2/Y V_GND 0.606f
C15134 FULL_COUNTER.COUNT_SUB_DFF4.Q V_GND 3.65f
C15135 sky130_fd_sc_hd__conb_1_0/HI V_GND 3.14f
C15136 sky130_fd_sc_hd__conb_1_3/HI V_GND 0.305f
C15137 sky130_fd_sc_hd__conb_1_4/HI V_GND 0.264f
C15138 sky130_fd_sc_hd__inv_1_3/Y V_GND 0.799f
C15139 sky130_fd_sc_hd__inv_1_0/Y V_GND 0.35f
C15140 FULL_COUNTER.COUNT_SUB_DFF2.Q V_GND 5.9f
C15141 sky130_fd_sc_hd__inv_16_40/Y V_GND 17.1f
C15142 sky130_fd_sc_hd__conb_1_5/HI V_GND 0.45f
C15143 sky130_fd_sc_hd__inv_1_14/Y V_GND 0.202f
C15144 sky130_fd_sc_hd__conb_1_10/HI V_GND 0.989f
C15145 sky130_fd_sc_hd__conb_1_9/HI V_GND 0.458f
C15146 sky130_fd_sc_hd__inv_1_9/Y V_GND 0.185f
C15147 sky130_fd_sc_hd__inv_1_13/Y V_GND 0.289f
C15148 sky130_fd_sc_hd__conb_1_14/HI V_GND 0.631f
C15149 sky130_fd_sc_hd__conb_1_7/HI V_GND 0.517f
C15150 sky130_fd_sc_hd__inv_1_7/Y V_GND 0.316f
C15151 RISING_COUNTER.COUNT_SUB_DFF15.Q V_GND 2.79f
C15152 sky130_fd_sc_hd__inv_1_21/Y V_GND 0.333f
C15153 sky130_fd_sc_hd__inv_1_69/Y V_GND 0.203f
C15154 sky130_fd_sc_hd__inv_16_4/Y V_GND 2.97f
C15155 sky130_fd_sc_hd__inv_4_0/A V_GND 0.907f
C15156 sky130_fd_sc_hd__inv_8_0/A V_GND 0.834f
C15157 sky130_fd_sc_hd__inv_16_9/A V_GND 1.74f
C15158 RISING_COUNTER.COUNT_SUB_DFF1.Q V_GND 5.84f
C15159 sky130_fd_sc_hd__inv_16_33/Y V_GND 1.61f
C15160 sky130_fd_sc_hd__conb_1_31/HI V_GND 0.379f
C15161 sky130_fd_sc_hd__inv_1_36/Y V_GND 0.576f
C15162 RISING_COUNTER.COUNT_SUB_DFF0.Q V_GND 6.28f
C15163 RISING_COUNTER.COUNT_SUB_DFF13.Q V_GND 1.52f
C15164 sky130_fd_sc_hd__nor2_1_0/Y V_GND 0.167f
C15165 sky130_fd_sc_hd__inv_2_0/A V_GND 0.933f
C15166 sky130_fd_sc_hd__nand2_8_8/A V_GND 0.684f
C15167 sky130_fd_sc_hd__inv_1_19/A V_GND 0.968f
C15168 sky130_fd_sc_hd__inv_1_46/A V_GND 2.97f
C15169 sky130_fd_sc_hd__inv_16_7/A V_GND 1.62f
C15170 sky130_fd_sc_hd__nand3_1_1/Y V_GND 1.01f
C15171 sky130_fd_sc_hd__inv_1_66/Y V_GND 1.44f
C15172 sky130_fd_sc_hd__inv_1_20/Y V_GND 1.14f
C15173 FALLING_COUNTER.COUNT_SUB_DFF13.Q V_GND 2.83f
C15174 sky130_fd_sc_hd__inv_1_53/A V_GND 0.952f
C15175 sky130_fd_sc_hd__conb_1_24/HI V_GND 0.832f
C15176 sky130_fd_sc_hd__inv_1_33/Y V_GND 0.526f
C15177 sky130_fd_sc_hd__inv_1_51/Y V_GND 0.757f
C15178 sky130_fd_sc_hd__inv_1_56/A V_GND 0.558f
C15179 sky130_fd_sc_hd__inv_1_53/Y V_GND 0.17f
C15180 sky130_fd_sc_hd__inv_1_23/Y V_GND 0.196f
C15181 FALLING_COUNTER.COUNT_SUB_DFF7.Q V_GND 1.68f
C15182 FALLING_COUNTER.COUNT_SUB_DFF2.Q V_GND 7.56f
C15183 FALLING_COUNTER.COUNT_SUB_DFF15.Q V_GND 1.98f
C15184 sky130_fd_sc_hd__inv_1_50/Y V_GND 0.215f
C15185 FALLING_COUNTER.COUNT_SUB_DFF12.Q V_GND 1.64f
C15186 sky130_fd_sc_hd__inv_1_61/Y V_GND 0.262f
C15187 sky130_fd_sc_hd__inv_1_63/Y V_GND 0.37f
C15188 sky130_fd_sc_hd__inv_1_62/Y V_GND 0.19f
C15189 sky130_fd_sc_hd__inv_16_19/Y V_GND 1.54f
C15190 sky130_fd_sc_hd__conb_1_47/HI V_GND 0.684f
C15191 sky130_fd_sc_hd__conb_1_46/HI V_GND 0.776f
C15192 sky130_fd_sc_hd__conb_1_41/HI V_GND 0.721f
C15193 FALLING_COUNTER.COUNT_SUB_DFF11.Q V_GND 1.7f
C15194 sky130_fd_sc_hd__conb_1_50/HI V_GND 0.421f
C15195 sky130_fd_sc_hd__inv_16_49/Y V_GND 7.32f
C15196 sky130_fd_sc_hd__inv_16_52/A V_GND 1.49f
C15197 sky130_fd_sc_hd__inv_1_12/Y V_GND 0.296f
C15198 sky130_fd_sc_hd__inv_1_32/Y V_GND 0.404f
C15199 sky130_fd_sc_hd__inv_1_18/A V_GND 1.14f
C15200 sky130_fd_sc_hd__inv_16_16/Y V_GND 1.61f
C15201 sky130_fd_sc_hd__dfbbn_1_5/Q_N V_GND 0.0166f
C15202 sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# V_GND 1.21e-19
C15203 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# V_GND 0.0118f
C15204 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# V_GND 0.14f
C15205 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# V_GND 1.77e-19
C15206 sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# V_GND 0.00102f
C15207 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# V_GND 2.96e-19
C15208 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# V_GND 0.0155f
C15209 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# V_GND 1.48e-19
C15210 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# V_GND 6.44e-19
C15211 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# V_GND 4.63e-19
C15212 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# V_GND 2.5e-19
C15213 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# V_GND 0.0255f
C15214 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# V_GND 0.126f
C15215 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# V_GND 0.404f
C15216 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# V_GND 0.254f
C15217 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# V_GND 0.125f
C15218 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# V_GND 0.246f
C15219 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# V_GND 0.283f
C15220 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# V_GND 0.547f
C15221 sky130_fd_sc_hd__inv_1_43/Y V_GND 0.336f
C15222 sky130_fd_sc_hd__nand2_8_1/a_27_47# V_GND 0.118f
C15223 sky130_fd_sc_hd__conb_1_12/HI V_GND 0.636f
C15224 sky130_fd_sc_hd__dfbbn_1_4/Q_N V_GND 0.0135f
C15225 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# V_GND 1.21e-19
C15226 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# V_GND 0.0116f
C15227 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# V_GND 0.139f
C15228 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# V_GND 4.81e-19
C15229 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# V_GND 0.00109f
C15230 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# V_GND -8.67e-19
C15231 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# V_GND 0.0156f
C15232 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# V_GND 2.66e-19
C15233 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# V_GND 0.00116f
C15234 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# V_GND 5.43e-19
C15235 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# V_GND 2.95e-19
C15236 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# V_GND 0.0184f
C15237 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# V_GND 0.127f
C15238 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# V_GND 0.401f
C15239 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# V_GND 0.231f
C15240 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# V_GND 0.119f
C15241 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# V_GND 0.248f
C15242 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# V_GND 0.278f
C15243 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# V_GND 0.356f
C15244 sky130_fd_sc_hd__nand2_8_9/A V_GND 0.735f
C15245 sky130_fd_sc_hd__nand2_8_4/Y V_GND 0.916f
C15246 sky130_fd_sc_hd__nand3_1_2/Y V_GND 0.956f
C15247 FALLING_COUNTER.COUNT_SUB_DFF10.Q V_GND 1.19f
C15248 sky130_fd_sc_hd__inv_1_60/Y V_GND 0.373f
C15249 sky130_fd_sc_hd__nand2_8_0/a_27_47# V_GND 0.131f
C15250 sky130_fd_sc_hd__conb_1_51/HI V_GND 1.06f
C15251 sky130_fd_sc_hd__conb_1_9/LO V_GND 0.169f
C15252 sky130_fd_sc_hd__fill_8_858/VPB V_GND 5.11f
C15253 sky130_fd_sc_hd__inv_1_11/Y V_GND 0.165f
C15254 sky130_fd_sc_hd__dfbbn_1_3/Q_N V_GND 0.01f
C15255 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# V_GND -1.67e-19
C15256 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# V_GND 0.00731f
C15257 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# V_GND 0.125f
C15258 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# V_GND 5.83e-19
C15259 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# V_GND -3.87e-19
C15260 sky130_fd_sc_hd__dfbbn_1_3/a_581_47# V_GND 7.87e-19
C15261 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# V_GND 0.0112f
C15262 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# V_GND 3.2e-19
C15263 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# V_GND 0.00142f
C15264 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# V_GND 6.31e-19
C15265 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# V_GND 4.04e-19
C15266 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# V_GND 0.0292f
C15267 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# V_GND 0.125f
C15268 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# V_GND 0.401f
C15269 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# V_GND 0.22f
C15270 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# V_GND 0.13f
C15271 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# V_GND 0.249f
C15272 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# V_GND 0.295f
C15273 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# V_GND 0.547f
C15274 sky130_fd_sc_hd__conb_1_39/HI V_GND 0.578f
C15275 sky130_fd_sc_hd__inv_1_47/A V_GND 1.24f
C15276 sky130_fd_sc_hd__inv_16_55/A V_GND 1.5f
C15277 sky130_fd_sc_hd__conb_1_8/LO V_GND 0.171f
C15278 sky130_fd_sc_hd__fill_8_848/VPB V_GND 5.11f
C15279 FALLING_COUNTER.COUNT_SUB_DFF14.Q V_GND 2.1f
C15280 sky130_fd_sc_hd__dfbbn_1_2/Q_N V_GND 0.0173f
C15281 sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# V_GND 5.2e-19
C15282 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# V_GND 0.0155f
C15283 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# V_GND 0.141f
C15284 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# V_GND 6.35e-19
C15285 sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# V_GND 0.00235f
C15286 sky130_fd_sc_hd__dfbbn_1_2/a_581_47# V_GND 7.48e-19
C15287 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# V_GND 0.0202f
C15288 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# V_GND 3.66e-19
C15289 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# V_GND 0.00192f
C15290 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# V_GND 0.00121f
C15291 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# V_GND 5.44e-19
C15292 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# V_GND 0.0283f
C15293 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# V_GND 0.135f
C15294 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# V_GND 0.414f
C15295 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# V_GND 0.274f
C15296 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# V_GND 0.134f
C15297 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# V_GND 0.257f
C15298 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# V_GND 0.292f
C15299 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# V_GND 0.547f
C15300 sky130_fd_sc_hd__inv_1_24/Y V_GND 1.28f
C15301 sky130_fd_sc_hd__nand2_1_5/a_113_47# V_GND 7.75e-20
C15302 sky130_fd_sc_hd__conb_1_35/HI V_GND 1.01f
C15303 sky130_fd_sc_hd__conb_1_7/LO V_GND 0.161f
C15304 sky130_fd_sc_hd__inv_1_65/Y V_GND 0.101f
C15305 sky130_fd_sc_hd__inv_16_48/Y V_GND 3.58f
C15306 sky130_fd_sc_hd__dfbbn_1_1/Q_N V_GND 0.0164f
C15307 sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# V_GND -1.67e-19
C15308 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# V_GND 0.00871f
C15309 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# V_GND 0.15f
C15310 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# V_GND 8.18e-19
C15311 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# V_GND -6.41e-19
C15312 sky130_fd_sc_hd__dfbbn_1_1/a_581_47# V_GND -6.92e-19
C15313 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# V_GND 0.0108f
C15314 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# V_GND 3.2e-19
C15315 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# V_GND 0.00142f
C15316 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# V_GND 6.31e-19
C15317 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# V_GND 3.4e-19
C15318 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# V_GND 0.0203f
C15319 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# V_GND 0.126f
C15320 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# V_GND 0.413f
C15321 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# V_GND 0.222f
C15322 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# V_GND 0.123f
C15323 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# V_GND 0.248f
C15324 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# V_GND 0.285f
C15325 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# V_GND 0.37f
C15326 sky130_fd_sc_hd__nand2_1_4/a_113_47# V_GND -5.45e-20
C15327 sky130_fd_sc_hd__conb_1_6/LO V_GND 0.168f
C15328 FULL_COUNTER.COUNT_SUB_DFF15.Q V_GND 4.73f
C15329 sky130_fd_sc_hd__dfbbn_1_0/Q_N V_GND 0.00585f
C15330 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# V_GND 2.1e-19
C15331 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# V_GND 0.00829f
C15332 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# V_GND 0.135f
C15333 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# V_GND 3.7e-19
C15334 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# V_GND 9.09e-19
C15335 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# V_GND 3.01e-19
C15336 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# V_GND 0.0148f
C15337 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# V_GND 3.24e-19
C15338 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# V_GND 0.00164f
C15339 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# V_GND 7.41e-19
C15340 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# V_GND 4.82e-19
C15341 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# V_GND 0.0244f
C15342 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# V_GND 0.127f
C15343 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# V_GND 0.396f
C15344 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# V_GND 0.222f
C15345 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# V_GND 0.125f
C15346 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# V_GND 0.247f
C15347 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# V_GND 0.282f
C15348 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# V_GND 0.507f
C15349 sky130_fd_sc_hd__nand2_1_3/Y V_GND 0.0488f
C15350 sky130_fd_sc_hd__nand2_1_3/a_113_47# V_GND -1.83e-19
C15351 sky130_fd_sc_hd__conb_1_5/LO V_GND 0.188f
C15352 sky130_fd_sc_hd__fill_8_854/VPB V_GND 5.13f
C15353 sky130_fd_sc_hd__inv_1_52/Y V_GND 0.0994f
C15354 sky130_fd_sc_hd__nand2_1_2/a_113_47# V_GND 1.94e-19
C15355 sky130_fd_sc_hd__conb_1_4/LO V_GND 0.165f
C15356 sky130_fd_sc_hd__nand2_1_1/a_113_47# V_GND -1.47e-19
C15357 sky130_fd_sc_hd__conb_1_3/LO V_GND 0.165f
C15358 sky130_fd_sc_hd__fill_8_852/VPB V_GND 5.11f
C15359 sky130_fd_sc_hd__conb_1_28/HI V_GND 0.26f
C15360 sky130_fd_sc_hd__inv_1_25/Y V_GND 0.307f
C15361 sky130_fd_sc_hd__nand2_1_0/a_113_47# V_GND 1.54e-19
C15362 sky130_fd_sc_hd__nand2_1_2/A V_GND 1.06f
C15363 sky130_fd_sc_hd__inv_1_42/Y V_GND 0.215f
C15364 sky130_fd_sc_hd__conb_1_19/LO V_GND 0.172f
C15365 sky130_fd_sc_hd__conb_1_2/LO V_GND 0.168f
C15366 sky130_fd_sc_hd__conb_1_18/LO V_GND 0.162f
C15367 sky130_fd_sc_hd__conb_1_29/LO V_GND 0.168f
C15368 sky130_fd_sc_hd__conb_1_1/LO V_GND 0.168f
C15369 sky130_fd_sc_hd__fill_4_189/VPB V_GND 5.04f
C15370 sky130_fd_sc_hd__fill_4_320/VPB V_GND 5.11f
C15371 sky130_fd_sc_hd__conb_1_39/LO V_GND 0.163f
C15372 sky130_fd_sc_hd__conb_1_17/LO V_GND 0.163f
C15373 sky130_fd_sc_hd__conb_1_28/LO V_GND 0.163f
C15374 sky130_fd_sc_hd__conb_1_0/LO V_GND 0.164f
C15375 sky130_fd_sc_hd__inv_16_5/A V_GND 1.51f
C15376 sky130_fd_sc_hd__conb_1_49/LO V_GND 0.172f
C15377 sky130_fd_sc_hd__conb_1_27/LO V_GND 0.169f
C15378 sky130_fd_sc_hd__conb_1_38/LO V_GND 0.171f
C15379 sky130_fd_sc_hd__conb_1_16/LO V_GND 0.166f
C15380 sky130_fd_sc_hd__fill_4_184/VPB V_GND 5.08f
C15381 sky130_fd_sc_hd__fill_4_194/VPB V_GND 5.09f
C15382 sky130_fd_sc_hd__inv_16_3/A V_GND 1.63f
C15383 sky130_fd_sc_hd__conb_1_48/LO V_GND 0.199f
C15384 sky130_fd_sc_hd__conb_1_26/LO V_GND 0.167f
C15385 sky130_fd_sc_hd__conb_1_37/LO V_GND 0.164f
C15386 sky130_fd_sc_hd__conb_1_15/LO V_GND 0.171f
C15387 RISING_COUNTER.COUNT_SUB_DFF11.Q V_GND 1.85f
C15388 sky130_fd_sc_hd__inv_16_27/Y V_GND 1.72f
C15389 sky130_fd_sc_hd__conb_1_47/LO V_GND 0.167f
C15390 sky130_fd_sc_hd__conb_1_25/LO V_GND 0.162f
C15391 sky130_fd_sc_hd__conb_1_36/LO V_GND 0.171f
C15392 sky130_fd_sc_hd__conb_1_14/LO V_GND 0.169f
C15393 sky130_fd_sc_hd__dfbbn_1_19/Q_N V_GND 0.0106f
C15394 sky130_fd_sc_hd__conb_1_20/HI V_GND 0.68f
C15395 sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# V_GND 2.51e-19
C15396 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# V_GND 0.0111f
C15397 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# V_GND 0.14f
C15398 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# V_GND 2.17e-19
C15399 sky130_fd_sc_hd__dfbbn_1_19/a_1159_47# V_GND 0.0011f
C15400 sky130_fd_sc_hd__dfbbn_1_19/a_581_47# V_GND 3.58e-19
C15401 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# V_GND 0.0152f
C15402 sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# V_GND 2.57e-19
C15403 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# V_GND 0.00157f
C15404 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# V_GND 7.07e-19
C15405 sky130_fd_sc_hd__dfbbn_1_19/a_557_413# V_GND 4.56e-19
C15406 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# V_GND 0.0246f
C15407 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# V_GND 0.124f
C15408 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# V_GND 0.396f
C15409 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# V_GND 0.209f
C15410 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# V_GND 0.126f
C15411 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# V_GND 0.248f
C15412 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# V_GND 0.283f
C15413 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# V_GND 0.539f
C15414 sky130_fd_sc_hd__inv_1_34/Y V_GND 0.331f
C15415 sky130_fd_sc_hd__conb_1_21/HI V_GND 0.848f
C15416 sky130_fd_sc_hd__conb_1_46/LO V_GND 0.169f
C15417 sky130_fd_sc_hd__conb_1_24/LO V_GND 0.167f
C15418 sky130_fd_sc_hd__conb_1_35/LO V_GND 0.162f
C15419 sky130_fd_sc_hd__conb_1_13/LO V_GND 0.171f
C15420 sky130_fd_sc_hd__inv_8_0/Y V_GND 1.61f
C15421 sky130_fd_sc_hd__dfbbn_1_29/Q_N V_GND 0.0124f
C15422 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# V_GND -4.04e-19
C15423 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# V_GND 0.00451f
C15424 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# V_GND 0.129f
C15425 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# V_GND 5.23e-19
C15426 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# V_GND -0.00126f
C15427 sky130_fd_sc_hd__dfbbn_1_29/a_581_47# V_GND 3.58e-19
C15428 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# V_GND 0.00859f
C15429 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# V_GND 2.55e-19
C15430 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# V_GND 0.00116f
C15431 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# V_GND 5.16e-19
C15432 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# V_GND 2.88e-19
C15433 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# V_GND 0.0245f
C15434 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# V_GND 0.117f
C15435 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# V_GND 0.393f
C15436 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# V_GND 0.205f
C15437 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# V_GND 0.122f
C15438 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# V_GND 0.242f
C15439 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# V_GND 0.281f
C15440 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# V_GND 0.498f
C15441 sky130_fd_sc_hd__dfbbn_1_18/Q_N V_GND 0.0139f
C15442 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# V_GND -2.77e-19
C15443 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# V_GND 0.00531f
C15444 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# V_GND 0.136f
C15445 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# V_GND 1.67e-19
C15446 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# V_GND -0.00114f
C15447 sky130_fd_sc_hd__dfbbn_1_18/a_581_47# V_GND -8.07e-19
C15448 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# V_GND 0.00953f
C15449 sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# V_GND 1.84e-19
C15450 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# V_GND 0.00107f
C15451 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# V_GND 4.8e-19
C15452 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# V_GND 2.82e-19
C15453 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# V_GND 0.0178f
C15454 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# V_GND 0.12f
C15455 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# V_GND 0.394f
C15456 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# V_GND 0.209f
C15457 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# V_GND 0.119f
C15458 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# V_GND 0.243f
C15459 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# V_GND 0.278f
C15460 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# V_GND 0.33f
C15461 RISING_COUNTER.COUNT_SUB_DFF9.Q V_GND 2.62f
C15462 sky130_fd_sc_hd__inv_1_23/A V_GND 1.02f
C15463 sky130_fd_sc_hd__inv_16_6/Y V_GND 1.55f
C15464 sky130_fd_sc_hd__conb_1_23/LO V_GND 0.17f
C15465 sky130_fd_sc_hd__conb_1_45/LO V_GND 0.165f
C15466 sky130_fd_sc_hd__conb_1_34/LO V_GND 0.162f
C15467 sky130_fd_sc_hd__conb_1_12/LO V_GND 0.171f
C15468 sky130_fd_sc_hd__inv_16_7/Y V_GND 1.66f
C15469 sky130_fd_sc_hd__inv_1_22/Y V_GND 0.919f
C15470 sky130_fd_sc_hd__dfbbn_1_39/Q_N V_GND 0.0142f
C15471 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# V_GND 2.48e-19
C15472 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# V_GND 0.0118f
C15473 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# V_GND 0.134f
C15474 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# V_GND 4.81e-19
C15475 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# V_GND 6.74e-19
C15476 sky130_fd_sc_hd__dfbbn_1_39/a_581_47# V_GND 3.54e-19
C15477 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# V_GND 0.0152f
C15478 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# V_GND 3.09e-19
C15479 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# V_GND 0.00158f
C15480 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# V_GND 7.12e-19
C15481 sky130_fd_sc_hd__dfbbn_1_39/a_557_413# V_GND 4.59e-19
C15482 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# V_GND 0.025f
C15483 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# V_GND 0.129f
C15484 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# V_GND 0.4f
C15485 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# V_GND 0.255f
C15486 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# V_GND 0.126f
C15487 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# V_GND 0.247f
C15488 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# V_GND 0.294f
C15489 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# V_GND 0.518f
C15490 sky130_fd_sc_hd__dfbbn_1_17/Q_N V_GND 0.00684f
C15491 sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# V_GND 2.11e-19
C15492 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# V_GND 0.0111f
C15493 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# V_GND 0.121f
C15494 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# V_GND 4.8e-19
C15495 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# V_GND 8.97e-19
C15496 sky130_fd_sc_hd__dfbbn_1_17/a_581_47# V_GND 3.29e-19
C15497 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# V_GND 0.0148f
C15498 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# V_GND 2.58e-19
C15499 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# V_GND 0.00157f
C15500 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# V_GND 7.09e-19
C15501 sky130_fd_sc_hd__dfbbn_1_17/a_557_413# V_GND 4.58e-19
C15502 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# V_GND 0.0243f
C15503 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# V_GND 0.138f
C15504 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# V_GND 0.405f
C15505 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# V_GND 0.211f
C15506 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# V_GND 0.125f
C15507 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# V_GND 0.247f
C15508 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# V_GND 0.284f
C15509 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# V_GND 0.519f
C15510 sky130_fd_sc_hd__dfbbn_1_28/Q_N V_GND 0.0185f
C15511 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# V_GND 1.52e-19
C15512 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# V_GND 0.0133f
C15513 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# V_GND 0.144f
C15514 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# V_GND 4.8e-19
C15515 sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# V_GND 0.00144f
C15516 sky130_fd_sc_hd__dfbbn_1_28/a_581_47# V_GND 4.66e-19
C15517 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# V_GND 0.0167f
C15518 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# V_GND 3.01e-19
C15519 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# V_GND 0.00148f
C15520 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# V_GND 6.71e-19
C15521 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# V_GND 4.48e-19
C15522 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# V_GND 0.0264f
C15523 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# V_GND 0.127f
C15524 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# V_GND 0.408f
C15525 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# V_GND 0.22f
C15526 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# V_GND 0.128f
C15527 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# V_GND 0.25f
C15528 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# V_GND 0.286f
C15529 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# V_GND 0.528f
C15530 sky130_fd_sc_hd__inv_1_55/Y V_GND 0.198f
C15531 sky130_fd_sc_hd__fill_4_182/VPB V_GND 5.1f
C15532 sky130_fd_sc_hd__fill_4_188/VPB V_GND 5.08f
C15533 sky130_fd_sc_hd__conb_1_44/LO V_GND 0.167f
C15534 sky130_fd_sc_hd__conb_1_33/LO V_GND 0.175f
C15535 sky130_fd_sc_hd__conb_1_22/LO V_GND 0.175f
C15536 sky130_fd_sc_hd__conb_1_11/LO V_GND 0.163f
C15537 sky130_fd_sc_hd__dfbbn_1_49/Q_N V_GND 0.0089f
C15538 sky130_fd_sc_hd__conb_1_45/HI V_GND 0.997f
C15539 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# V_GND 2.51e-19
C15540 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# V_GND 0.0118f
C15541 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# V_GND 0.121f
C15542 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# V_GND 3.29e-19
C15543 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# V_GND 0.00109f
C15544 sky130_fd_sc_hd__dfbbn_1_49/a_581_47# V_GND -8.5e-19
C15545 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# V_GND 0.0151f
C15546 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# V_GND 1.89e-19
C15547 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# V_GND 0.00116f
C15548 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# V_GND 5.16e-19
C15549 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# V_GND 2.88e-19
C15550 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# V_GND 0.0172f
C15551 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# V_GND 0.127f
C15552 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# V_GND 0.401f
C15553 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# V_GND 0.251f
C15554 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# V_GND 0.118f
C15555 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# V_GND 0.261f
C15556 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# V_GND 0.276f
C15557 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# V_GND 0.347f
C15558 sky130_fd_sc_hd__dfbbn_1_38/Q_N V_GND 0.00735f
C15559 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# V_GND -3.18e-19
C15560 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# V_GND 0.00443f
C15561 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# V_GND 0.135f
C15562 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# V_GND 5.23e-19
C15563 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# V_GND -0.00126f
C15564 sky130_fd_sc_hd__dfbbn_1_38/a_581_47# V_GND 3.57e-19
C15565 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# V_GND 0.00955f
C15566 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# V_GND 3.09e-19
C15567 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# V_GND 0.00158f
C15568 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# V_GND 7.12e-19
C15569 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# V_GND 4.59e-19
C15570 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# V_GND 0.025f
C15571 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# V_GND 0.118f
C15572 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# V_GND 0.391f
C15573 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# V_GND 0.205f
C15574 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# V_GND 0.134f
C15575 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# V_GND 0.244f
C15576 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# V_GND 0.281f
C15577 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# V_GND 0.518f
C15578 sky130_fd_sc_hd__dfbbn_1_27/Q_N V_GND 0.0144f
C15579 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# V_GND 2.51e-19
C15580 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# V_GND 0.0107f
C15581 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# V_GND 0.137f
C15582 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# V_GND 5.12e-19
C15583 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# V_GND 0.00109f
C15584 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# V_GND 3.57e-19
C15585 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# V_GND 0.0152f
C15586 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# V_GND 2.53e-19
C15587 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# V_GND 0.00152f
C15588 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# V_GND 6.9e-19
C15589 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# V_GND 4.48e-19
C15590 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# V_GND 0.0245f
C15591 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# V_GND 0.124f
C15592 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# V_GND 0.4f
C15593 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# V_GND 0.212f
C15594 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# V_GND 0.126f
C15595 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# V_GND 0.248f
C15596 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# V_GND 0.283f
C15597 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# V_GND 0.507f
C15598 sky130_fd_sc_hd__dfbbn_1_16/Q_N V_GND 0.00623f
C15599 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# V_GND 2.45e-19
C15600 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# V_GND 0.00656f
C15601 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# V_GND 0.122f
C15602 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# V_GND 2.5e-19
C15603 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# V_GND 0.00104f
C15604 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# V_GND 3.49e-19
C15605 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# V_GND 0.015f
C15606 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# V_GND 4.09e-19
C15607 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# V_GND 0.00209f
C15608 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# V_GND 9.44e-19
C15609 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# V_GND 6.09e-19
C15610 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# V_GND 0.0262f
C15611 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# V_GND 0.125f
C15612 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# V_GND 0.395f
C15613 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# V_GND 0.213f
C15614 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# V_GND 0.127f
C15615 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# V_GND 0.25f
C15616 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# V_GND 0.295f
C15617 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# V_GND 0.515f
C15618 RISING_COUNTER.COUNT_SUB_DFF7.Q V_GND 6.02f
C15619 sky130_fd_sc_hd__conb_1_18/HI V_GND 0.644f
C15620 sky130_fd_sc_hd__inv_1_52/A V_GND 0.961f
C15621 sky130_fd_sc_hd__nand3_1_2/a_193_47# V_GND -8.64e-19
C15622 sky130_fd_sc_hd__nand3_1_2/a_109_47# V_GND -4.72e-19
C15623 sky130_fd_sc_hd__conb_1_43/LO V_GND 0.167f
C15624 sky130_fd_sc_hd__conb_1_32/LO V_GND 0.164f
C15625 sky130_fd_sc_hd__conb_1_21/LO V_GND 0.17f
C15626 sky130_fd_sc_hd__conb_1_10/LO V_GND 0.167f
C15627 sky130_fd_sc_hd__inv_1_8/Y V_GND 0.363f
C15628 sky130_fd_sc_hd__dfbbn_1_26/Q_N V_GND 0.0105f
C15629 sky130_fd_sc_hd__conb_1_25/HI V_GND 0.643f
C15630 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# V_GND 1.2e-19
C15631 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# V_GND 0.0127f
C15632 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# V_GND 0.135f
C15633 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# V_GND 2.18e-19
C15634 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# V_GND 0.00108f
C15635 sky130_fd_sc_hd__dfbbn_1_26/a_581_47# V_GND 3.54e-19
C15636 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# V_GND 0.0151f
C15637 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# V_GND 2.6e-19
C15638 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# V_GND 0.00158f
C15639 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# V_GND 7.12e-19
C15640 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# V_GND 4.59e-19
C15641 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# V_GND 0.0238f
C15642 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# V_GND 0.126f
C15643 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# V_GND 0.409f
C15644 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# V_GND 0.21f
C15645 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# V_GND 0.125f
C15646 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# V_GND 0.248f
C15647 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# V_GND 0.281f
C15648 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# V_GND 0.539f
C15649 sky130_fd_sc_hd__dfbbn_1_48/Q_N V_GND 0.0174f
C15650 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# V_GND -3.2e-19
C15651 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# V_GND 0.0043f
C15652 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# V_GND 0.142f
C15653 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# V_GND 2.6e-19
C15654 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# V_GND -0.00132f
C15655 sky130_fd_sc_hd__dfbbn_1_48/a_581_47# V_GND -8.52e-19
C15656 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# V_GND 0.0086f
C15657 sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# V_GND 3.09e-19
C15658 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# V_GND 0.00108f
C15659 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# V_GND 7.12e-19
C15660 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# V_GND 4.59e-19
C15661 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# V_GND 0.018f
C15662 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# V_GND 0.118f
C15663 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# V_GND 0.4f
C15664 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# V_GND 0.208f
C15665 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# V_GND 0.117f
C15666 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# V_GND 0.242f
C15667 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# V_GND 0.276f
C15668 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# V_GND 0.346f
C15669 sky130_fd_sc_hd__dfbbn_1_37/Q_N V_GND 0.00702f
C15670 sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# V_GND -3.48e-19
C15671 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# V_GND 0.00409f
C15672 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# V_GND 0.121f
C15673 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# V_GND 5.21e-19
C15674 sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# V_GND -0.00142f
C15675 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# V_GND -8.65e-19
C15676 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# V_GND 0.008f
C15677 sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# V_GND 3.08e-19
C15678 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# V_GND 0.00157f
C15679 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# V_GND 6.98e-19
C15680 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# V_GND 4.58e-19
C15681 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# V_GND 0.018f
C15682 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# V_GND 0.119f
C15683 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# V_GND 0.391f
C15684 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# V_GND 0.202f
C15685 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# V_GND 0.116f
C15686 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# V_GND 0.242f
C15687 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# V_GND 0.275f
C15688 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# V_GND 0.323f
C15689 sky130_fd_sc_hd__dfbbn_1_15/Q_N V_GND 0.0122f
C15690 sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# V_GND 2.5e-19
C15691 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# V_GND 0.0118f
C15692 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# V_GND 0.129f
C15693 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# V_GND 4.16e-19
C15694 sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# V_GND 0.00109f
C15695 sky130_fd_sc_hd__dfbbn_1_15/a_581_47# V_GND 3.57e-19
C15696 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# V_GND 0.0154f
C15697 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# V_GND 2.19e-19
C15698 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# V_GND 0.00139f
C15699 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# V_GND 6.26e-19
C15700 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# V_GND 3.95e-19
C15701 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# V_GND 0.0246f
C15702 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# V_GND 0.124f
C15703 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# V_GND 0.397f
C15704 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# V_GND 0.214f
C15705 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# V_GND 0.126f
C15706 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# V_GND 0.247f
C15707 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# V_GND 0.282f
C15708 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# V_GND 0.532f
C15709 FALLING_COUNTER.COUNT_SUB_DFF8.Q V_GND 1.35f
C15710 sky130_fd_sc_hd__inv_16_42/Y V_GND 12.2f
C15711 sky130_fd_sc_hd__conb_1_43/HI V_GND 0.356f
C15712 sky130_fd_sc_hd__nand3_1_1/a_193_47# V_GND -6.18e-19
C15713 sky130_fd_sc_hd__nand3_1_1/a_109_47# V_GND -5.01e-20
C15714 sky130_fd_sc_hd__inv_16_26/A V_GND 1.45f
C15715 sky130_fd_sc_hd__conb_1_42/LO V_GND 0.18f
C15716 sky130_fd_sc_hd__conb_1_20/LO V_GND 0.17f
C15717 sky130_fd_sc_hd__conb_1_31/LO V_GND 0.173f
C15718 sky130_fd_sc_hd__inv_1_4/Y V_GND 0.528f
C15719 sky130_fd_sc_hd__dfbbn_1_25/Q_N V_GND 0.00735f
C15720 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# V_GND -3.18e-19
C15721 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# V_GND 0.00406f
C15722 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# V_GND 0.124f
C15723 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# V_GND 4.81e-19
C15724 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# V_GND -0.00142f
C15725 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# V_GND 3.57e-19
C15726 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# V_GND 0.00864f
C15727 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# V_GND 2.59e-19
C15728 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# V_GND 0.00108f
C15729 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# V_GND 7.12e-19
C15730 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# V_GND 4.59e-19
C15731 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# V_GND 0.0238f
C15732 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# V_GND 0.117f
C15733 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# V_GND 0.389f
C15734 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# V_GND 0.201f
C15735 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# V_GND 0.121f
C15736 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# V_GND 0.242f
C15737 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# V_GND 0.278f
C15738 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# V_GND 0.515f
C15739 sky130_fd_sc_hd__dfbbn_1_47/Q_N V_GND 0.00737f
C15740 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# V_GND 1.21e-19
C15741 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# V_GND 0.00832f
C15742 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# V_GND 0.124f
C15743 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# V_GND 5.12e-19
C15744 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# V_GND 0.00109f
C15745 sky130_fd_sc_hd__dfbbn_1_47/a_581_47# V_GND 3.57e-19
C15746 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# V_GND 0.0152f
C15747 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# V_GND 3.02e-19
C15748 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# V_GND 0.00152f
C15749 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# V_GND 6.97e-19
C15750 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# V_GND 4.48e-19
C15751 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# V_GND 0.0246f
C15752 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# V_GND 0.125f
C15753 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# V_GND 0.393f
C15754 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# V_GND 0.205f
C15755 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# V_GND 0.126f
C15756 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# V_GND 0.248f
C15757 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# V_GND 0.282f
C15758 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# V_GND 0.508f
C15759 sky130_fd_sc_hd__dfbbn_1_36/Q_N V_GND 0.00804f
C15760 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# V_GND 4.24e-19
C15761 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# V_GND 0.0103f
C15762 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# V_GND 0.123f
C15763 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# V_GND 4.81e-19
C15764 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# V_GND 0.00255f
C15765 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# V_GND -7.49e-19
C15766 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# V_GND 0.0169f
C15767 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# V_GND 2.47e-19
C15768 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# V_GND 0.00224f
C15769 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# V_GND 7.58e-19
C15770 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# V_GND 4.19e-19
C15771 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# V_GND 0.0188f
C15772 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# V_GND 0.131f
C15773 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# V_GND 0.398f
C15774 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# V_GND 0.227f
C15775 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# V_GND 0.121f
C15776 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# V_GND 0.252f
C15777 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# V_GND 0.282f
C15778 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# V_GND 0.354f
C15779 sky130_fd_sc_hd__dfbbn_1_14/Q_N V_GND 0.0065f
C15780 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# V_GND -3.19e-19
C15781 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# V_GND 0.00382f
C15782 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# V_GND 0.125f
C15783 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# V_GND 2.6e-19
C15784 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# V_GND -0.00126f
C15785 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# V_GND 3.55e-19
C15786 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# V_GND 0.00841f
C15787 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# V_GND 3.09e-19
C15788 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# V_GND 0.00158f
C15789 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# V_GND 7.05e-19
C15790 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# V_GND 4.59e-19
C15791 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# V_GND 0.0245f
C15792 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# V_GND 0.118f
C15793 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# V_GND 0.4f
C15794 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# V_GND 0.202f
C15795 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# V_GND 0.122f
C15796 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# V_GND 0.243f
C15797 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# V_GND 0.28f
C15798 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# V_GND 0.516f
C15799 sky130_fd_sc_hd__fill_4_215/VPB V_GND 5.09f
C15800 sky130_fd_sc_hd__nand3_1_0/a_193_47# V_GND -7.36e-19
C15801 sky130_fd_sc_hd__nand3_1_0/a_109_47# V_GND -5.05e-19
C15802 sky130_fd_sc_hd__conb_1_41/LO V_GND 0.173f
C15803 sky130_fd_sc_hd__conb_1_30/LO V_GND 0.163f
C15804 sky130_fd_sc_hd__dfbbn_1_46/Q_N V_GND 0.00613f
C15805 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# V_GND -4.04e-19
C15806 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# V_GND 0.00609f
C15807 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# V_GND 0.122f
C15808 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# V_GND 5.23e-19
C15809 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# V_GND -0.00131f
C15810 sky130_fd_sc_hd__dfbbn_1_46/a_581_47# V_GND -8.5e-19
C15811 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# V_GND 0.00852f
C15812 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# V_GND 3.04e-19
C15813 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# V_GND 0.00108f
C15814 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# V_GND 7.12e-19
C15815 sky130_fd_sc_hd__dfbbn_1_46/a_557_413# V_GND 4.59e-19
C15816 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# V_GND 0.0176f
C15817 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# V_GND 0.12f
C15818 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# V_GND 0.389f
C15819 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# V_GND 0.203f
C15820 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# V_GND 0.117f
C15821 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# V_GND 0.242f
C15822 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# V_GND 0.275f
C15823 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# V_GND 0.316f
C15824 sky130_fd_sc_hd__dfbbn_1_35/Q_N V_GND 0.00584f
C15825 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# V_GND -4.07e-19
C15826 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# V_GND 0.00386f
C15827 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# V_GND 0.122f
C15828 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# V_GND 4.8e-19
C15829 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# V_GND -0.00172f
C15830 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# V_GND -8.88e-19
C15831 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# V_GND 0.00733f
C15832 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# V_GND 2.58e-19
C15833 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# V_GND 0.00157f
C15834 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# V_GND 7.09e-19
C15835 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# V_GND 4.58e-19
C15836 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# V_GND 0.0175f
C15837 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# V_GND 0.117f
C15838 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# V_GND 0.387f
C15839 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# V_GND 0.201f
C15840 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# V_GND 0.115f
C15841 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# V_GND 0.24f
C15842 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# V_GND 0.274f
C15843 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# V_GND 0.347f
C15844 sky130_fd_sc_hd__dfbbn_1_24/Q_N V_GND 0.0161f
C15845 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# V_GND -3.2e-19
C15846 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# V_GND 0.00392f
C15847 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# V_GND 0.14f
C15848 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# V_GND 2.6e-19
C15849 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# V_GND -0.00132f
C15850 sky130_fd_sc_hd__dfbbn_1_24/a_581_47# V_GND -8.52e-19
C15851 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# V_GND 0.00846f
C15852 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# V_GND 3.09e-19
C15853 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# V_GND 0.00108f
C15854 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# V_GND 7.12e-19
C15855 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# V_GND 4.59e-19
C15856 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# V_GND 0.018f
C15857 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# V_GND 0.118f
C15858 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# V_GND 0.396f
C15859 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# V_GND 0.203f
C15860 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# V_GND 0.116f
C15861 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# V_GND 0.242f
C15862 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# V_GND 0.275f
C15863 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# V_GND 0.315f
C15864 sky130_fd_sc_hd__dfbbn_1_13/Q_N V_GND 0.00766f
C15865 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# V_GND 2.45e-19
C15866 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# V_GND 0.0107f
C15867 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# V_GND 0.12f
C15868 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# V_GND 4.91e-19
C15869 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# V_GND 0.00104f
C15870 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# V_GND 3.49e-19
C15871 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# V_GND 0.0151f
C15872 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# V_GND 2.14e-19
C15873 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# V_GND 0.00154f
C15874 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# V_GND 6.84e-19
C15875 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# V_GND 3.82e-19
C15876 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# V_GND 0.0253f
C15877 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# V_GND 0.126f
C15878 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# V_GND 0.4f
C15879 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# V_GND 0.215f
C15880 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# V_GND 0.126f
C15881 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# V_GND 0.249f
C15882 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# V_GND 0.292f
C15883 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# V_GND 0.524f
C15884 sky130_fd_sc_hd__conb_1_33/HI V_GND 0.323f
C15885 sky130_fd_sc_hd__conb_1_44/HI V_GND 0.664f
C15886 RISING_COUNTER.COUNT_SUB_DFF12.Q V_GND 2.77f
C15887 sky130_fd_sc_hd__inv_1_68/Y V_GND 0.345f
C15888 sky130_fd_sc_hd__inv_16_32/A V_GND 1.77f
C15889 sky130_fd_sc_hd__conb_1_51/LO V_GND 0.163f
C15890 sky130_fd_sc_hd__conb_1_40/LO V_GND 0.173f
C15891 sky130_fd_sc_hd__dfbbn_1_45/Q_N V_GND 0.0145f
C15892 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# V_GND 3.64e-19
C15893 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# V_GND 0.0129f
C15894 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# V_GND 0.144f
C15895 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# V_GND 6.28e-19
C15896 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# V_GND 0.00136f
C15897 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# V_GND 5.4e-19
C15898 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# V_GND 0.0164f
C15899 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# V_GND 4.15e-19
C15900 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# V_GND 0.00205f
C15901 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# V_GND 9.29e-19
C15902 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# V_GND 6.17e-19
C15903 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# V_GND 0.0269f
C15904 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# V_GND 0.132f
C15905 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# V_GND 0.407f
C15906 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# V_GND 0.265f
C15907 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# V_GND 0.131f
C15908 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# V_GND 0.25f
C15909 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# V_GND 0.29f
C15910 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# V_GND 0.54f
C15911 sky130_fd_sc_hd__dfbbn_1_34/Q_N V_GND 0.0185f
C15912 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# V_GND 3.64e-19
C15913 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# V_GND 0.0137f
C15914 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# V_GND 0.143f
C15915 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# V_GND 4.66e-19
C15916 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# V_GND 0.00185f
C15917 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# V_GND -7.81e-19
C15918 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# V_GND 0.0169f
C15919 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# V_GND 2.28e-19
C15920 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# V_GND 0.00192f
C15921 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# V_GND 6.67e-19
C15922 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# V_GND 3.89e-19
C15923 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# V_GND 0.0192f
C15924 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# V_GND 0.131f
C15925 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# V_GND 0.411f
C15926 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# V_GND 0.265f
C15927 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# V_GND 0.122f
C15928 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# V_GND 0.25f
C15929 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# V_GND 0.28f
C15930 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# V_GND 0.361f
C15931 sky130_fd_sc_hd__dfbbn_1_23/Q_N V_GND 0.0107f
C15932 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# V_GND -3.18e-19
C15933 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# V_GND 0.00676f
C15934 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# V_GND 0.128f
C15935 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# V_GND 3.71e-19
C15936 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# V_GND -0.00137f
C15937 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# V_GND -8.97e-19
C15938 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# V_GND 0.0083f
C15939 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# V_GND 1.89e-19
C15940 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# V_GND 0.00116f
C15941 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# V_GND 5.16e-19
C15942 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# V_GND 2.19e-19
C15943 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# V_GND 0.0175f
C15944 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# V_GND 0.119f
C15945 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# V_GND 0.392f
C15946 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# V_GND 0.209f
C15947 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# V_GND 0.116f
C15948 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# V_GND 0.241f
C15949 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# V_GND 0.274f
C15950 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# V_GND 0.313f
C15951 sky130_fd_sc_hd__dfbbn_1_12/Q_N V_GND 0.0174f
C15952 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# V_GND 2.5e-19
C15953 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# V_GND 0.0118f
C15954 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# V_GND 0.142f
C15955 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# V_GND 5.23e-19
C15956 sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# V_GND 9.3e-19
C15957 sky130_fd_sc_hd__dfbbn_1_12/a_581_47# V_GND 3.57e-19
C15958 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# V_GND 0.0153f
C15959 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# V_GND 2.59e-19
C15960 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# V_GND 0.00108f
C15961 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# V_GND 7.12e-19
C15962 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# V_GND 4.59e-19
C15963 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# V_GND 0.025f
C15964 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# V_GND 0.125f
C15965 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# V_GND 0.408f
C15966 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# V_GND 0.214f
C15967 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# V_GND 0.126f
C15968 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# V_GND 0.247f
C15969 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# V_GND 0.282f
C15970 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# V_GND 0.509f
C15971 sky130_fd_sc_hd__conb_1_48/HI V_GND 0.443f
C15972 sky130_fd_sc_hd__conb_1_34/HI V_GND 0.243f
C15973 FALLING_COUNTER.COUNT_SUB_DFF1.Q V_GND 6.18f
C15974 sky130_fd_sc_hd__inv_1_54/Y V_GND 0.257f
C15975 sky130_fd_sc_hd__inv_1_67/Y V_GND 1.01f
C15976 sky130_fd_sc_hd__nand2_8_9/Y V_GND 0.744f
C15977 sky130_fd_sc_hd__conb_1_50/LO V_GND 0.163f
C15978 sky130_fd_sc_hd__dfbbn_1_44/Q_N V_GND 0.014f
C15979 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# V_GND -3.48e-19
C15980 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# V_GND 0.00403f
C15981 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# V_GND 0.133f
C15982 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# V_GND 4.8e-19
C15983 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# V_GND -0.00146f
C15984 sky130_fd_sc_hd__dfbbn_1_44/a_581_47# V_GND 3.29e-19
C15985 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# V_GND 0.00823f
C15986 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# V_GND 2.58e-19
C15987 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# V_GND 0.00108f
C15988 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# V_GND 7.09e-19
C15989 sky130_fd_sc_hd__dfbbn_1_44/a_557_413# V_GND 4.58e-19
C15990 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# V_GND 0.0243f
C15991 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# V_GND 0.118f
C15992 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# V_GND 0.394f
C15993 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# V_GND 0.203f
C15994 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# V_GND 0.123f
C15995 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# V_GND 0.242f
C15996 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# V_GND 0.281f
C15997 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# V_GND 0.526f
C15998 sky130_fd_sc_hd__dfbbn_1_22/Q_N V_GND 0.0162f
C15999 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# V_GND 2.49e-19
C16000 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# V_GND 0.0113f
C16001 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# V_GND 0.14f
C16002 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# V_GND 5.6e-19
C16003 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# V_GND 8.29e-19
C16004 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# V_GND -8.51e-19
C16005 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# V_GND 0.0153f
C16006 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# V_GND 2.82e-19
C16007 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# V_GND 0.00121f
C16008 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# V_GND 7.84e-19
C16009 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# V_GND 5.18e-19
C16010 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# V_GND 0.0169f
C16011 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# V_GND 0.127f
C16012 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# V_GND 0.403f
C16013 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# V_GND 0.255f
C16014 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# V_GND 0.118f
C16015 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# V_GND 0.247f
C16016 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# V_GND 0.274f
C16017 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# V_GND 0.344f
C16018 sky130_fd_sc_hd__dfbbn_1_33/Q_N V_GND 0.0157f
C16019 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# V_GND -3.48e-19
C16020 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# V_GND 0.00403f
C16021 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# V_GND 0.138f
C16022 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# V_GND 3.28e-19
C16023 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# V_GND -0.00142f
C16024 sky130_fd_sc_hd__dfbbn_1_33/a_581_47# V_GND -8.65e-19
C16025 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# V_GND 0.00818f
C16026 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# V_GND 1.73e-19
C16027 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# V_GND 0.00157f
C16028 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# V_GND 7.09e-19
C16029 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# V_GND 4.58e-19
C16030 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# V_GND 0.0177f
C16031 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# V_GND 0.117f
C16032 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# V_GND 0.396f
C16033 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# V_GND 0.202f
C16034 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# V_GND 0.117f
C16035 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# V_GND 0.243f
C16036 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# V_GND 0.274f
C16037 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# V_GND 0.314f
C16038 sky130_fd_sc_hd__dfbbn_1_11/Q_N V_GND 0.00849f
C16039 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# V_GND -3.21e-19
C16040 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# V_GND 0.00439f
C16041 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# V_GND 0.127f
C16042 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# V_GND 4.91e-19
C16043 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# V_GND -0.0013f
C16044 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# V_GND -8.54e-19
C16045 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# V_GND 0.00856f
C16046 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# V_GND 2.5e-19
C16047 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# V_GND 0.00154f
C16048 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# V_GND 6.84e-19
C16049 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# V_GND 3.82e-19
C16050 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# V_GND 0.0187f
C16051 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# V_GND 0.12f
C16052 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# V_GND 0.397f
C16053 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# V_GND 0.212f
C16054 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# V_GND 0.119f
C16055 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# V_GND 0.244f
C16056 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# V_GND 0.288f
C16057 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# V_GND 0.337f
C16058 sky130_fd_sc_hd__inv_1_37/Y V_GND 0.312f
C16059 sky130_fd_sc_hd__conb_1_42/HI V_GND 0.673f
C16060 sky130_fd_sc_hd__fill_8_958/VPB V_GND 5.11f
C16061 sky130_fd_sc_hd__dfbbn_1_43/Q_N V_GND 0.00708f
C16062 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# V_GND -3.18e-19
C16063 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# V_GND 0.00443f
C16064 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# V_GND 0.12f
C16065 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# V_GND 3.71e-19
C16066 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# V_GND -0.00126f
C16067 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# V_GND -8.5e-19
C16068 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# V_GND 0.00838f
C16069 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# V_GND 1.62e-19
C16070 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# V_GND 0.00116f
C16071 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# V_GND 5.16e-19
C16072 sky130_fd_sc_hd__dfbbn_1_43/a_557_413# V_GND 2.88e-19
C16073 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# V_GND 0.0176f
C16074 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# V_GND 0.12f
C16075 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# V_GND 0.398f
C16076 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# V_GND 0.202f
C16077 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# V_GND 0.116f
C16078 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# V_GND 0.242f
C16079 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# V_GND 0.277f
C16080 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# V_GND 0.344f
C16081 sky130_fd_sc_hd__dfbbn_1_21/Q_N V_GND 0.0175f
C16082 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# V_GND 1.2e-19
C16083 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# V_GND 0.0118f
C16084 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# V_GND 0.14f
C16085 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# V_GND 5.88e-19
C16086 sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# V_GND 8.67e-19
C16087 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# V_GND 2.26e-19
C16088 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# V_GND 0.015f
C16089 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# V_GND 3.41e-19
C16090 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# V_GND 0.00171f
C16091 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# V_GND 7.84e-19
C16092 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# V_GND 3.94e-19
C16093 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# V_GND 0.0247f
C16094 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# V_GND 0.126f
C16095 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# V_GND 0.409f
C16096 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# V_GND 0.214f
C16097 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# V_GND 0.126f
C16098 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# V_GND 0.247f
C16099 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# V_GND 0.285f
C16100 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# V_GND 0.505f
C16101 sky130_fd_sc_hd__dfbbn_1_32/Q_N V_GND 0.0121f
C16102 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# V_GND 3.24e-19
C16103 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# V_GND 0.0125f
C16104 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# V_GND 0.141f
C16105 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# V_GND 4.53e-19
C16106 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# V_GND 0.00144f
C16107 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# V_GND 6.21e-19
C16108 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# V_GND 0.0167f
C16109 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# V_GND 3.01e-19
C16110 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# V_GND 0.00148f
C16111 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# V_GND 0.00118f
C16112 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# V_GND 7.89e-19
C16113 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# V_GND 0.0269f
C16114 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# V_GND 0.127f
C16115 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# V_GND 0.411f
C16116 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# V_GND 0.214f
C16117 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# V_GND 0.131f
C16118 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# V_GND 0.252f
C16119 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# V_GND 0.288f
C16120 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# V_GND 0.559f
C16121 sky130_fd_sc_hd__dfbbn_1_10/Q_N V_GND 0.0113f
C16122 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# V_GND -4.04e-19
C16123 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# V_GND 0.00442f
C16124 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# V_GND 0.127f
C16125 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# V_GND 5.23e-19
C16126 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# V_GND -0.00135f
C16127 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# V_GND -8.51e-19
C16128 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# V_GND 0.00847f
C16129 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# V_GND 3.04e-19
C16130 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# V_GND 0.00158f
C16131 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# V_GND 7.12e-19
C16132 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# V_GND 4.59e-19
C16133 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# V_GND 0.0177f
C16134 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# V_GND 0.117f
C16135 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# V_GND 0.39f
C16136 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# V_GND 0.202f
C16137 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# V_GND 0.116f
C16138 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# V_GND 0.241f
C16139 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# V_GND 0.273f
C16140 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# V_GND 0.313f
C16141 sky130_fd_sc_hd__dfbbn_1_42/Q_N V_GND 0.0168f
C16142 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# V_GND -3.18e-19
C16143 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# V_GND 0.00535f
C16144 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# V_GND 0.14f
C16145 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# V_GND 3.71e-19
C16146 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# V_GND -0.00131f
C16147 sky130_fd_sc_hd__dfbbn_1_42/a_581_47# V_GND -8.5e-19
C16148 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# V_GND 0.00852f
C16149 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# V_GND 1.89e-19
C16150 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# V_GND 7.71e-19
C16151 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# V_GND 5.16e-19
C16152 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# V_GND 2.88e-19
C16153 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# V_GND 0.0189f
C16154 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# V_GND 0.129f
C16155 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# V_GND 0.401f
C16156 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# V_GND 0.207f
C16157 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# V_GND 0.117f
C16158 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# V_GND 0.242f
C16159 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# V_GND 0.286f
C16160 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# V_GND 0.314f
C16161 sky130_fd_sc_hd__dfbbn_1_31/Q_N V_GND 0.00703f
C16162 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# V_GND -3.48e-19
C16163 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# V_GND 0.00361f
C16164 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# V_GND 0.122f
C16165 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# V_GND 2.59e-19
C16166 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# V_GND -0.00142f
C16167 sky130_fd_sc_hd__dfbbn_1_31/a_581_47# V_GND 3.29e-19
C16168 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# V_GND 0.00817f
C16169 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# V_GND 3.08e-19
C16170 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# V_GND 0.00157f
C16171 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# V_GND 7.09e-19
C16172 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# V_GND 3.46e-19
C16173 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# V_GND 0.0246f
C16174 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# V_GND 0.117f
C16175 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# V_GND 0.388f
C16176 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# V_GND 0.202f
C16177 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# V_GND 0.121f
C16178 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# V_GND 0.242f
C16179 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# V_GND 0.281f
C16180 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# V_GND 0.518f
C16181 sky130_fd_sc_hd__dfbbn_1_20/Q_N V_GND 0.0172f
C16182 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# V_GND 3.24e-19
C16183 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# V_GND 0.0133f
C16184 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# V_GND 0.144f
C16185 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# V_GND 4.53e-19
C16186 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# V_GND 0.00119f
C16187 sky130_fd_sc_hd__dfbbn_1_20/a_581_47# V_GND 4.66e-19
C16188 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# V_GND 0.0178f
C16189 sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# V_GND 3.01e-19
C16190 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# V_GND 0.00148f
C16191 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# V_GND 6.71e-19
C16192 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# V_GND 4.48e-19
C16193 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# V_GND 0.026f
C16194 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# V_GND 0.13f
C16195 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# V_GND 0.408f
C16196 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# V_GND 0.275f
C16197 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# V_GND 0.129f
C16198 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# V_GND 0.252f
C16199 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# V_GND 0.288f
C16200 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# V_GND 0.565f
C16201 sky130_fd_sc_hd__fill_8_932/VPB V_GND 5.11f
C16202 sky130_fd_sc_hd__dfbbn_1_41/Q_N V_GND 0.0174f
C16203 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# V_GND 2.48e-19
C16204 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# V_GND 0.0118f
C16205 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# V_GND 0.138f
C16206 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# V_GND 5.23e-19
C16207 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# V_GND 0.00108f
C16208 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# V_GND 3.54e-19
C16209 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# V_GND 0.0152f
C16210 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# V_GND 2.59e-19
C16211 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# V_GND 0.00158f
C16212 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# V_GND 7e-19
C16213 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# V_GND 4.59e-19
C16214 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# V_GND 0.025f
C16215 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# V_GND 0.127f
C16216 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# V_GND 0.406f
C16217 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# V_GND 0.256f
C16218 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# V_GND 0.125f
C16219 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# V_GND 0.247f
C16220 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# V_GND 0.282f
C16221 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# V_GND 0.508f
C16222 sky130_fd_sc_hd__dfbbn_1_30/Q_N V_GND 0.0116f
C16223 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# V_GND -3.48e-19
C16224 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# V_GND 0.00417f
C16225 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# V_GND 0.147f
C16226 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# V_GND 5.21e-19
C16227 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# V_GND -0.00146f
C16228 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# V_GND -8.65e-19
C16229 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# V_GND 0.00824f
C16230 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# V_GND 3.08e-19
C16231 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# V_GND 0.00108f
C16232 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# V_GND 7.09e-19
C16233 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# V_GND 4.58e-19
C16234 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# V_GND 0.017f
C16235 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# V_GND 0.117f
C16236 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# V_GND 0.398f
C16237 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# V_GND 0.203f
C16238 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# V_GND 0.117f
C16239 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# V_GND 0.243f
C16240 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# V_GND 0.273f
C16241 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# V_GND 0.315f
C16242 sky130_fd_sc_hd__inv_1_65/A V_GND 0.931f
C16243 sky130_fd_sc_hd__conb_1_13/HI V_GND 0.371f
C16244 sky130_fd_sc_hd__dfbbn_1_51/Q_N V_GND 0.0174f
C16245 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# V_GND -3.2e-19
C16246 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# V_GND 0.00445f
C16247 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# V_GND 0.139f
C16248 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# V_GND 5.23e-19
C16249 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# V_GND -0.00127f
C16250 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# V_GND -8.52e-19
C16251 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# V_GND 0.0086f
C16252 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# V_GND 2.59e-19
C16253 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# V_GND 0.00158f
C16254 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# V_GND 7.12e-19
C16255 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# V_GND 4.59e-19
C16256 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# V_GND 0.0177f
C16257 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# V_GND 0.119f
C16258 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# V_GND 0.401f
C16259 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# V_GND 0.202f
C16260 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# V_GND 0.117f
C16261 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# V_GND 0.243f
C16262 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# V_GND 0.275f
C16263 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# V_GND 0.316f
C16264 sky130_fd_sc_hd__dfbbn_1_40/Q_N V_GND 0.00737f
C16265 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# V_GND 2.48e-19
C16266 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# V_GND 0.0118f
C16267 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# V_GND 0.123f
C16268 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# V_GND 4.81e-19
C16269 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# V_GND 9.19e-19
C16270 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# V_GND 3.54e-19
C16271 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# V_GND 0.0153f
C16272 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# V_GND 3.09e-19
C16273 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# V_GND 0.00108f
C16274 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# V_GND 7.12e-19
C16275 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# V_GND 4.59e-19
C16276 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# V_GND 0.025f
C16277 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# V_GND 0.127f
C16278 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# V_GND 0.398f
C16279 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# V_GND 0.254f
C16280 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# V_GND 0.126f
C16281 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# V_GND 0.247f
C16282 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# V_GND 0.283f
C16283 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# V_GND 0.542f
C16284 sky130_fd_sc_hd__conb_1_22/HI V_GND 0.74f
C16285 sky130_fd_sc_hd__inv_16_20/A V_GND 2.06f
C16286 sky130_fd_sc_hd__dfbbn_1_50/Q_N V_GND 0.00831f
C16287 sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# V_GND 3.24e-19
C16288 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# V_GND 0.013f
C16289 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# V_GND 0.125f
C16290 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# V_GND 4.8e-19
C16291 sky130_fd_sc_hd__dfbbn_1_50/a_1159_47# V_GND 0.00118f
C16292 sky130_fd_sc_hd__dfbbn_1_50/a_581_47# V_GND 4.66e-19
C16293 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# V_GND 0.0164f
C16294 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# V_GND 3.01e-19
C16295 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# V_GND 0.00148f
C16296 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# V_GND 6.71e-19
C16297 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# V_GND 4.48e-19
C16298 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# V_GND 0.0263f
C16299 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# V_GND 0.13f
C16300 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# V_GND 0.413f
C16301 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# V_GND 0.233f
C16302 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# V_GND 0.128f
C16303 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# V_GND 0.249f
C16304 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# V_GND 0.285f
C16305 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# V_GND 0.557f
C16306 sky130_fd_sc_hd__inv_16_23/Y V_GND 1.67f
C16307 sky130_fd_sc_hd__conb_1_1/HI V_GND 0.623f
C16308 sky130_fd_sc_hd__inv_1_15/Y V_GND 0.299f
C16309 RISING_COUNTER.COUNT_SUB_DFF14.Q V_GND 2.03f
C16310 sky130_fd_sc_hd__inv_16_44/Y V_GND 2.73f
C16311 sky130_fd_sc_hd__fill_8_951/VPB V_GND 5.11f
C16312 sky130_fd_sc_hd__fill_8_927/VPB V_GND 5.12f
C16313 sky130_fd_sc_hd__nand2_8_9/a_27_47# V_GND 0.0969f
C16314 sky130_fd_sc_hd__conb_1_49/HI V_GND 0.435f
C16315 sky130_fd_sc_hd__inv_16_45/A V_GND 2.36f
C16316 sky130_fd_sc_hd__inv_16_26/Y V_GND 1.44f
C16317 sky130_fd_sc_hd__nand2_8_8/a_27_47# V_GND 0.135f
C16318 sky130_fd_sc_hd__nand3_1_0/Y V_GND 1.48f
C16319 sky130_fd_sc_hd__inv_16_31/Y V_GND 1.48f
C16320 sky130_fd_sc_hd__nor2_1_0/a_109_297# V_GND -7.26e-19
C16321 sky130_fd_sc_hd__conb_1_36/HI V_GND 0.288f
C16322 sky130_fd_sc_hd__nand2_8_7/a_27_47# V_GND 0.114f
C16323 FULL_COUNTER.COUNT_SUB_DFF19.Q V_GND 4.79f
C16324 sky130_fd_sc_hd__inv_16_6/A V_GND 13.4f
C16325 sky130_fd_sc_hd__nand2_8_6/a_27_47# V_GND 0.0281f
C16326 sky130_fd_sc_hd__inv_1_18/Y V_GND 0.101f
C16327 sky130_fd_sc_hd__dfbbn_1_9/Q_N V_GND 0.0144f
C16328 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# V_GND 1.21e-19
C16329 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# V_GND 0.0118f
C16330 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# V_GND 0.134f
C16331 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# V_GND 5.23e-19
C16332 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# V_GND 8.74e-19
C16333 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# V_GND 2.96e-19
C16334 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# V_GND 0.0155f
C16335 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# V_GND 3.04e-19
C16336 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# V_GND 0.00158f
C16337 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# V_GND 7.48e-19
C16338 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# V_GND 4.67e-19
C16339 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# V_GND 0.0263f
C16340 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# V_GND 0.127f
C16341 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# V_GND 0.401f
C16342 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# V_GND 0.255f
C16343 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# V_GND 0.127f
C16344 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# V_GND 0.248f
C16345 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# V_GND 0.285f
C16346 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# V_GND 0.549f
C16347 sky130_fd_sc_hd__inv_1_57/Y V_GND 0.355f
C16348 sky130_fd_sc_hd__nand2_8_5/a_27_47# V_GND 0.139f
C16349 sky130_fd_sc_hd__inv_1_6/Y V_GND 0.282f
C16350 V_SENSE V_GND 0.399p
C16351 sky130_fd_sc_hd__inv_16_23/A V_GND 1.73f
C16352 sky130_fd_sc_hd__inv_16_50/Y V_GND 5.16f
C16353 sky130_fd_sc_hd__dfbbn_1_8/Q_N V_GND 0.00698f
C16354 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# V_GND -3.19e-19
C16355 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# V_GND 0.00443f
C16356 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# V_GND 0.122f
C16357 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# V_GND 5.23e-19
C16358 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# V_GND -0.00135f
C16359 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# V_GND 3.55e-19
C16360 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# V_GND 0.00847f
C16361 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# V_GND 2.59e-19
C16362 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# V_GND 0.00158f
C16363 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# V_GND 7.12e-19
C16364 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# V_GND 4.59e-19
C16365 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# V_GND 0.0246f
C16366 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# V_GND 0.118f
C16367 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# V_GND 0.389f
C16368 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# V_GND 0.203f
C16369 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# V_GND 0.121f
C16370 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# V_GND 0.242f
C16371 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# V_GND 0.28f
C16372 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# V_GND 0.485f
C16373 sky130_fd_sc_hd__fill_8_949/VPB V_GND 5.12f
C16374 sky130_fd_sc_hd__nand2_8_4/a_27_47# V_GND 0.13f
C16375 sky130_fd_sc_hd__inv_1_16/Y V_GND 0.253f
C16376 sky130_fd_sc_hd__inv_16_44/A V_GND 2.4f
C16377 sky130_fd_sc_hd__inv_16_14/Y V_GND 1.68f
C16378 sky130_fd_sc_hd__dfbbn_1_7/Q_N V_GND 0.0181f
C16379 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# V_GND -3.19e-19
C16380 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# V_GND 0.00477f
C16381 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# V_GND 0.143f
C16382 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# V_GND 6.89e-19
C16383 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# V_GND -0.00138f
C16384 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# V_GND 3.55e-19
C16385 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# V_GND 0.00841f
C16386 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# V_GND 2.59e-19
C16387 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# V_GND 0.00158f
C16388 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# V_GND 7.12e-19
C16389 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# V_GND 4.59e-19
C16390 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# V_GND 0.0244f
C16391 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# V_GND 0.12f
C16392 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# V_GND 0.415f
C16393 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# V_GND 0.202f
C16394 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# V_GND 0.122f
C16395 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# V_GND 0.246f
C16396 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# V_GND 0.284f
C16397 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# V_GND 0.496f
C16398 RISING_COUNTER.COUNT_SUB_DFF2.Q V_GND 6.54f
C16399 sky130_fd_sc_hd__nand2_8_3/a_27_47# V_GND 0.116f
C16400 sky130_fd_sc_hd__inv_1_5/Y V_GND 0.243f
C16401 FULL_COUNTER.COUNT_SUB_DFF3.Q V_GND 2.92f
C16402 sky130_fd_sc_hd__dfbbn_1_6/Q_N V_GND 0.013f
C16403 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# V_GND 2.45e-19
C16404 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# V_GND 0.0117f
C16405 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# V_GND 0.136f
C16406 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# V_GND 4.91e-19
C16407 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# V_GND 8.58e-19
C16408 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# V_GND -8.54e-19
C16409 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# V_GND 0.0151f
C16410 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# V_GND 2.5e-19
C16411 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# V_GND 0.00154f
C16412 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# V_GND 6.84e-19
C16413 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# V_GND 3.82e-19
C16414 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# V_GND 0.0183f
C16415 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# V_GND 0.129f
C16416 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# V_GND 0.407f
C16417 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# V_GND 0.264f
C16418 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# V_GND 0.12f
C16419 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# V_GND 0.249f
C16420 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# V_GND 0.285f
C16421 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# V_GND 0.353f
C16422 sky130_fd_sc_hd__nand2_8_2/a_27_47# V_GND 0.139f
.ends
