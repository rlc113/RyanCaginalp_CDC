VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO transmission_gate
  CLASS Core ;
  FOREIGN transmission_gate ;
  ORIGIN 0 0 ;
  SIZE 3.22 BY 2.72 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN O
    ANTENNADIFFAREA 0.451000 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.600 2.220 2.100 ;
        RECT 1.980 0.940 2.190 1.600 ;
        RECT 1.870 0.640 2.220 0.940 ;
        RECT 2.410 0.640 2.800 0.910 ;
        RECT 1.870 0.440 2.800 0.640 ;
    END
  END O
  PIN G
    ANTENNAGATEAREA 0.082500 ;
    PORT
      LAYER li1 ;
        RECT 2.510 1.080 2.900 1.530 ;
    END
  END G
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.185 1.310 3.415 2.910 ;
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN GN
    ANTENNAGATEAREA 0.082500 ;
    PORT
      LAYER li1 ;
        RECT 2.460 2.110 2.850 2.560 ;
    END
  END GN
  OBS
      LAYER li1 ;
        RECT 0.700 2.080 1.110 2.910 ;
        RECT 0.660 1.630 1.110 2.080 ;
        RECT 0.750 1.420 1.110 1.630 ;
        RECT 1.310 1.600 1.660 2.100 ;
        RECT 1.370 1.420 1.600 1.600 ;
        RECT 0.560 1.170 1.600 1.420 ;
        RECT 1.370 0.940 1.600 1.170 ;
        RECT 0.660 0.470 1.110 0.920 ;
        RECT 0.710 -0.200 1.090 0.470 ;
        RECT 1.310 0.440 1.660 0.940 ;
      LAYER mcon ;
        RECT 0.780 2.520 1.070 2.860 ;
        RECT 0.770 -0.130 1.040 0.180 ;
  END
END transmission_gate
END LIBRARY

