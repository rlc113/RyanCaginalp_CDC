* NGSPICE file created from CDC.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_8 VNB VPB VGND VPWR A Y B a_27_47#
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B A 0.051f
C1 B VGND 0.108f
C2 B VPWR 0.118f
C3 B a_27_47# 0.369f
C4 B Y 0.413f
C5 VPB A 0.247f
C6 VPB VGND 0.0101f
C7 VPB VPWR 0.157f
C8 VPB a_27_47# 0.00278f
C9 VPB Y 0.0366f
C10 A VGND 0.0645f
C11 A VPWR 0.129f
C12 A a_27_47# 0.0695f
C13 VPB B 0.248f
C14 VPWR VGND 0.149f
C15 A Y 0.644f
C16 VGND a_27_47# 0.947f
C17 VPWR a_27_47# 0.0392f
C18 Y VGND 0.0559f
C19 VPWR Y 1.49f
C20 Y a_27_47# 0.337f
C21 VGND VNB 0.797f
C22 Y VNB 0.0446f
C23 VPWR VNB 0.753f
C24 A VNB 0.746f
C25 B VNB 0.758f
C26 VPB VNB 1.49f
C27 a_27_47# VNB 0.083f
.ends

.subckt sky130_fd_sc_hd__decap_4 VNB VPB VGND VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VPB VGND 0.116f
C1 VPB VPWR 0.0787f
C2 VGND VPWR 0.546f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__dfbbn_1 VNB VPB VGND VPWR Q Q_N RESET_B SET_B D CLK_N a_2136_47#
+ a_791_47# a_647_21# a_891_329# a_1363_47# a_557_413# a_941_21# a_1415_315# a_473_413#
+ a_193_47# a_381_47# a_1112_329# a_1555_47# a_581_47# a_1340_413# a_1159_47# a_1256_413#
+ a_1672_329# a_27_47#
X0 a_791_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0974 pd=0.97 as=0.0882 ps=0.84 w=0.42 l=0.15
X1 a_1555_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.03 as=0.0703 ps=0.755 w=0.42 l=0.15
X2 VPWR RESET_B a_941_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.17 ps=1.81 w=0.64 l=0.15
X3 a_1415_315# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.132 pd=1.22 as=0.0956 ps=0.875 w=0.42 l=0.15
X4 a_791_47# a_941_21# a_647_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5 VGND a_1415_315# a_1363_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.066 ps=0.745 w=0.42 l=0.15
X6 a_1340_413# a_27_47# a_1256_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0787 pd=0.795 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_473_413# a_193_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0675 pd=0.735 as=0.066 ps=0.745 w=0.36 l=0.15
X10 a_1555_47# a_941_21# a_1415_315# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VPWR a_1415_315# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_1256_413# a_193_47# a_1112_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X13 a_581_47# a_27_47# a_473_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0675 ps=0.735 w=0.36 l=0.15
X14 a_647_21# a_473_413# a_791_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X15 a_647_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X16 VPWR a_941_21# a_891_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X17 a_557_413# a_193_47# a_473_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X20 a_473_413# a_27_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0651 ps=0.73 w=0.42 l=0.15
X21 a_891_329# a_473_413# a_647_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X22 Q_N a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X23 VGND RESET_B a_941_21# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X24 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X25 VPWR a_647_21# a_557_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X26 a_1112_329# a_647_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X27 VGND a_647_21# a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X28 VGND a_1415_315# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 VPWR a_941_21# a_1672_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X31 VPWR a_1415_315# a_1340_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0956 pd=0.875 as=0.0787 ps=0.795 w=0.42 l=0.15
X32 a_1363_47# a_193_47# a_1256_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0486 ps=0.63 w=0.36 l=0.15
X33 Q_N a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X35 a_1159_47# a_647_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.116 pd=1.09 as=0.166 ps=1.8 w=0.64 l=0.15
X36 a_1672_329# a_1256_413# a_1415_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.132 ps=1.22 w=0.84 l=0.15
X37 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X38 a_1256_413# a_27_47# a_1159_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0486 pd=0.63 as=0.116 ps=1.09 w=0.36 l=0.15
X39 a_1415_315# a_1256_413# a_1555_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.109 ps=1.03 w=0.64 l=0.15
C0 a_27_47# a_791_47# 0.00134f
C1 a_473_413# VPWR 0.108f
C2 a_941_21# D 1.12e-19
C3 a_27_47# D 0.11f
C4 Q a_2136_47# 0.0721f
C5 VPB D 0.0817f
C6 a_381_47# D 0.148f
C7 a_647_21# a_891_329# 0.0104f
C8 a_1256_413# VPWR 0.12f
C9 a_193_47# Q 5.52e-20
C10 SET_B a_1363_47# 7.87e-19
C11 a_647_21# a_473_413# 0.206f
C12 a_473_413# VGND 0.147f
C13 a_941_21# VPWR 0.197f
C14 a_27_47# a_581_47# 0.00206f
C15 VPWR a_27_47# 0.146f
C16 VPWR VPB 0.255f
C17 a_381_47# a_581_47# 3.81e-19
C18 VPWR a_381_47# 0.0894f
C19 a_647_21# a_1256_413# 0.00189f
C20 a_193_47# a_1112_329# 0.00907f
C21 a_1256_413# a_1159_47# 0.00386f
C22 a_1256_413# VGND 0.127f
C23 a_647_21# a_941_21# 0.199f
C24 a_647_21# a_27_47# 0.15f
C25 a_941_21# a_1159_47# 3.73e-19
C26 a_1415_315# VPWR 0.315f
C27 a_473_413# RESET_B 7.48e-21
C28 a_941_21# VGND 0.134f
C29 a_27_47# a_1159_47# 0.00272f
C30 VGND a_27_47# 0.292f
C31 a_647_21# VPB 0.141f
C32 a_1555_47# a_1363_47# 4.19e-20
C33 VPWR CLK_N 0.0196f
C34 VGND VPB 0.0151f
C35 a_647_21# a_381_47# 8.07e-20
C36 VGND a_381_47# 0.0775f
C37 a_557_413# VPWR 0.0042f
C38 a_473_413# SET_B 0.14f
C39 a_1256_413# RESET_B 4.43e-20
C40 a_941_21# a_1672_329# 0.0016f
C41 a_941_21# RESET_B 0.105f
C42 RESET_B a_27_47# 2.12e-19
C43 a_1415_315# VGND 0.0797f
C44 RESET_B VPB 0.0476f
C45 VGND CLK_N 0.0196f
C46 VPWR D 0.0153f
C47 a_647_21# a_557_413# 6.69e-20
C48 a_193_47# a_891_329# 0.00276f
C49 a_1256_413# SET_B 0.177f
C50 RESET_B a_381_47# 3.34e-21
C51 a_193_47# a_473_413# 0.15f
C52 a_941_21# SET_B 0.096f
C53 SET_B a_27_47# 0.309f
C54 a_1256_413# Q_N 1e-20
C55 SET_B VPB 0.147f
C56 a_941_21# Q_N 0.0054f
C57 a_1415_315# a_1672_329# 0.00869f
C58 a_1415_315# RESET_B 0.0851f
C59 a_647_21# a_791_47# 0.0697f
C60 a_941_21# a_2136_47# 5.84e-19
C61 Q_N a_27_47# 4.78e-20
C62 a_27_47# a_2136_47# 1.76e-19
C63 a_791_47# a_1159_47# 3.34e-19
C64 VGND a_791_47# 0.164f
C65 a_2136_47# VPB 0.0467f
C66 Q_N VPB 0.0102f
C67 VGND D 0.0134f
C68 a_193_47# a_1256_413# 0.0334f
C69 a_193_47# a_941_21# 0.126f
C70 a_193_47# a_27_47# 0.798f
C71 a_1415_315# SET_B 0.141f
C72 a_1256_413# a_1555_47# 0.0256f
C73 a_193_47# VPB 0.198f
C74 a_193_47# a_381_47# 0.189f
C75 a_1415_315# a_2136_47# 0.0967f
C76 a_941_21# a_1555_47# 0.0526f
C77 a_1415_315# Q_N 0.121f
C78 a_647_21# VPWR 0.16f
C79 a_941_21# Q 1.7e-19
C80 Q a_27_47# 2.71e-20
C81 VGND a_581_47# 0.0017f
C82 VPWR a_1159_47# 6.2e-19
C83 VPWR VGND 0.0801f
C84 a_1555_47# VPB 8.96e-20
C85 Q VPB 0.0123f
C86 a_193_47# a_1415_315# 0.0494f
C87 a_1256_413# a_1112_329# 0.00412f
C88 a_193_47# CLK_N 7.87e-19
C89 a_1256_413# a_1363_47# 0.00707f
C90 SET_B a_791_47# 0.03f
C91 a_193_47# a_557_413# 0.0018f
C92 a_941_21# a_1112_329# 0.00652f
C93 a_1112_329# a_27_47# 1.09e-19
C94 a_647_21# a_1159_47# 9.75e-19
C95 a_941_21# a_1363_47# 1.96e-20
C96 a_647_21# VGND 0.053f
C97 a_1415_315# a_1555_47# 0.0383f
C98 a_1415_315# Q 0.00311f
C99 VPWR a_1672_329# 0.00438f
C100 VPWR RESET_B 0.0099f
C101 VGND a_1159_47# 0.0108f
C102 a_1256_413# a_1340_413# 0.00857f
C103 a_193_47# a_791_47# 6.04e-20
C104 a_193_47# D 0.0986f
C105 SET_B VPWR 0.0255f
C106 a_941_21# a_1340_413# 9.41e-19
C107 a_1340_413# a_27_47# 2.13e-19
C108 a_647_21# RESET_B 6.51e-21
C109 VPWR a_2136_47# 0.139f
C110 VPWR Q_N 0.0614f
C111 VGND RESET_B 0.0282f
C112 a_941_21# a_891_329# 1.21e-20
C113 a_891_329# a_27_47# 2.46e-19
C114 a_647_21# SET_B 0.175f
C115 a_193_47# VPWR 0.443f
C116 SET_B a_1159_47# 0.00459f
C117 SET_B VGND 0.311f
C118 a_473_413# a_941_21# 0.0633f
C119 a_473_413# a_27_47# 0.159f
C120 a_473_413# VPB 0.0627f
C121 a_791_47# a_1363_47# 2.46e-21
C122 VGND Q_N 0.0862f
C123 VGND a_2136_47# 0.114f
C124 VPWR a_1555_47# 1.3e-19
C125 VPWR Q 0.0992f
C126 a_473_413# a_381_47# 0.0369f
C127 a_193_47# a_647_21# 0.117f
C128 a_941_21# a_1256_413# 0.13f
C129 a_1256_413# a_27_47# 0.14f
C130 a_193_47# a_1159_47# 2.14e-20
C131 a_193_47# VGND 0.0661f
C132 a_1256_413# VPB 0.0597f
C133 SET_B RESET_B 0.00229f
C134 a_473_413# a_1415_315# 4.59e-22
C135 a_941_21# a_27_47# 0.14f
C136 a_941_21# VPB 0.142f
C137 a_1112_329# VPWR 0.0164f
C138 a_27_47# VPB 0.224f
C139 Q_N a_1672_329# 2.1e-20
C140 RESET_B a_2136_47# 4.99e-19
C141 RESET_B Q_N 0.0017f
C142 VGND a_1555_47# 0.157f
C143 VGND Q 0.0643f
C144 a_941_21# a_381_47# 3.79e-20
C145 a_381_47# a_27_47# 0.0456f
C146 a_473_413# a_557_413# 0.00972f
C147 a_381_47# VPB 0.0197f
C148 a_1415_315# a_1256_413# 0.207f
C149 a_193_47# a_1672_329# 7.17e-20
C150 a_193_47# RESET_B 6.8e-20
C151 SET_B a_2136_47# 3.22e-19
C152 SET_B Q_N 3.72e-19
C153 a_1415_315# a_27_47# 0.0321f
C154 a_941_21# a_1415_315# 0.267f
C155 a_647_21# a_1112_329# 9.46e-19
C156 a_473_413# a_791_47# 0.025f
C157 a_1340_413# VPWR 0.00281f
C158 a_1112_329# VGND 3.84e-19
C159 a_941_21# CLK_N 5.45e-20
C160 a_473_413# D 1.43e-19
C161 a_27_47# CLK_N 0.212f
C162 a_1415_315# VPB 0.242f
C163 Q_N a_2136_47# 0.175f
C164 VGND a_1363_47# 0.00192f
C165 RESET_B a_1555_47# 3.78e-20
C166 RESET_B Q 6.25e-20
C167 VPB CLK_N 0.0706f
C168 a_557_413# a_27_47# 4.45e-20
C169 a_193_47# SET_B 0.0123f
C170 a_557_413# a_381_47# 8.99e-19
C171 a_193_47# a_2136_47# 1.03e-19
C172 a_1256_413# a_791_47# 0.00316f
C173 a_193_47# Q_N 1.07e-19
C174 a_891_329# VPWR 0.00984f
C175 SET_B a_1555_47# 0.0131f
C176 SET_B Q 1.24e-19
C177 a_941_21# a_791_47# 0.00926f
C178 a_473_413# a_581_47# 0.00807f
C179 Q VNB 0.0945f
C180 Q_N VNB 0.0135f
C181 RESET_B VNB 0.133f
C182 VGND VNB 1.3f
C183 VPWR VNB 1.05f
C184 SET_B VNB 0.264f
C185 D VNB 0.125f
C186 CLK_N VNB 0.197f
C187 VPB VNB 2.38f
C188 a_1555_47# VNB 0.00871f
C189 a_2136_47# VNB 0.133f
C190 a_791_47# VNB 0.0125f
C191 a_381_47# VNB 0.0218f
C192 a_1256_413# VNB 0.12f
C193 a_1415_315# VNB 0.394f
C194 a_941_21# VNB 0.245f
C195 a_473_413# VNB 0.119f
C196 a_647_21# VNB 0.24f
C197 a_193_47# VNB 0.27f
C198 a_27_47# VNB 0.492f
.ends

.subckt sky130_fd_sc_hd__inv_1 VNB VPB VGND VPWR A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
C0 Y VGND 0.0998f
C1 VPB A 0.0451f
C2 VPB VPWR 0.0545f
C3 A VPWR 0.037f
C4 VPB Y 0.0177f
C5 VPB VGND 0.00948f
C6 A Y 0.0476f
C7 A VGND 0.04f
C8 VPWR Y 0.128f
C9 VPWR VGND 0.0338f
C10 VGND VNB 0.251f
C11 Y VNB 0.0961f
C12 VPWR VNB 0.219f
C13 A VNB 0.167f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nor2_1 VNB VPB VGND VPWR A B Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 A Y 0.0471f
C1 VPWR a_109_297# 0.00638f
C2 VGND a_109_297# 0.00128f
C3 VGND VPWR 0.0314f
C4 VPB VPWR 0.0449f
C5 B VPWR 0.0148f
C6 VGND VPB 0.00456f
C7 A VPWR 0.0528f
C8 Y a_109_297# 0.0113f
C9 VGND B 0.0451f
C10 Y VPWR 0.0995f
C11 VPB B 0.0367f
C12 VGND A 0.0486f
C13 VPB A 0.0415f
C14 VGND Y 0.154f
C15 B A 0.0584f
C16 VPB Y 0.0139f
C17 B Y 0.0877f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__inv_2 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 A Y 0.0894f
C1 VPB VGND 0.00649f
C2 VGND VPWR 0.0423f
C3 A VGND 0.0638f
C4 Y VGND 0.155f
C5 VPB VPWR 0.0521f
C6 VPB A 0.0742f
C7 A VPWR 0.0631f
C8 VPB Y 0.0061f
C9 Y VPWR 0.209f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt transmission_gate G VPWR VGND O GN
X0 O G VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.226 pd=1.92 as=0.226 ps=1.92 w=0.55 l=0.15
X1 O GN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.226 pd=1.92 as=0.226 ps=1.92 w=0.55 l=0.15
C0 VPWR GN 0.231f
C1 VPWR G 0.0852f
C2 VPWR O 0.145f
C3 GN G 0.0448f
C4 GN O 0.0144f
C5 O G 0.0806f
C6 G VGND 0.207f
C7 O VGND 0.14f
C8 GN VGND 0.0973f
C9 VPWR VGND 1.14f
.ends

.subckt sky130_fd_sc_hd__conb_1 VNB VPB VGND VPWR LO HI
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
C0 VPB LO 0.134f
C1 VPWR HI 0.0726f
C2 VGND HI 0.207f
C3 VGND VPWR 0.0317f
C4 LO HI 0.0683f
C5 LO VPWR 0.241f
C6 LO VGND 0.0605f
C7 VPB HI 0.00473f
C8 VPB VPWR 0.158f
C9 VPB VGND 0.00479f
C10 VGND VNB 0.406f
C11 LO VNB 0.166f
C12 HI VNB 0.25f
C13 VPWR VNB 0.297f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nand3_1 VNB VPB VGND VPWR A B Y C a_193_47# a_109_47#
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 C B 0.051f
C1 VPWR Y 0.317f
C2 VPWR VGND 0.0416f
C3 Y VPB 0.0166f
C4 Y a_193_47# 0.0117f
C5 Y C 0.0724f
C6 VGND VPB 0.00519f
C7 VPWR a_109_47# 2.94e-19
C8 VGND a_193_47# 0.00142f
C9 Y B 0.149f
C10 VPWR A 0.0186f
C11 VGND C 0.0415f
C12 VGND B 0.0116f
C13 VPB A 0.0368f
C14 B a_109_47# 4.42e-19
C15 VPWR VPB 0.0506f
C16 B A 0.0823f
C17 VPWR a_193_47# 5.03e-19
C18 Y VGND 0.181f
C19 VPWR C 0.0414f
C20 Y a_109_47# 0.0108f
C21 VPWR B 0.017f
C22 VPB C 0.0373f
C23 Y A 0.0909f
C24 VGND a_109_47# 9.04e-19
C25 VPB B 0.0268f
C26 a_193_47# B 0.00347f
C27 VGND A 0.01f
C28 VGND VNB 0.263f
C29 Y VNB 0.0816f
C30 VPWR VNB 0.247f
C31 A VNB 0.143f
C32 B VNB 0.0976f
C33 C VNB 0.157f
C34 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__nand2_1 VNB VPB VGND VPWR A Y B a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 VPB VGND 0.0044f
C1 VPB A 0.0379f
C2 B Y 0.0481f
C3 A VGND 0.00949f
C4 VPB Y 0.00618f
C5 Y VGND 0.139f
C6 A Y 0.0855f
C7 a_113_47# VGND 0.0019f
C8 a_113_47# Y 0.00937f
C9 VPWR B 0.0478f
C10 VPB VPWR 0.0509f
C11 VPWR VGND 0.0322f
C12 A VPWR 0.0444f
C13 VPWR Y 0.211f
C14 a_113_47# VPWR 1.78e-19
C15 VPB B 0.0391f
C16 B VGND 0.0544f
C17 A B 0.051f
C18 VGND VNB 0.232f
C19 Y VNB 0.0557f
C20 VPWR VNB 0.245f
C21 A VNB 0.143f
C22 B VNB 0.146f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__inv_16 VNB VPB VGND VPWR Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 Y VGND 1.06f
C1 A VPWR 0.28f
C2 VPB A 0.526f
C3 A Y 1.43f
C4 A VGND 0.266f
C5 VPB VPWR 0.159f
C6 VPWR Y 1.47f
C7 VPB Y 0.0305f
C8 VPWR VGND 0.161f
C9 VPB VGND 0.0132f
C10 VGND VNB 0.865f
C11 Y VNB 0.0551f
C12 VPWR VNB 0.737f
C13 A VNB 1.55f
C14 VPB VNB 1.49f
.ends

.subckt CDC CLOCK_GEN.SR_Op.Q FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF10.Q
+ FULL_COUNTER.COUNT_SUB_DFF11.Q FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF13.Q
+ FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF16.Q
+ FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF18.Q FULL_COUNTER.COUNT_SUB_DFF19.Q
+ FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF3.Q
+ FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF6.Q
+ FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF9.Q
+ RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF11.Q
+ RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF14.Q
+ RISING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF2.Q
+ RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF4.Q RISING_COUNTER.COUNT_SUB_DFF5.Q
+ RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF8.Q
+ RISING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q
+ FALLING_COUNTER.COUNT_SUB_DFF13.Q FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF15.Q
+ V_GND V_HIGH V_SENSE FALLING_COUNTER.COUNT_SUB_DFF0.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q
+ FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q
+ FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_DFF6.Q
+ FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q
+ Reset V_LOW
Xsky130_fd_sc_hd__nand2_8_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_8_2/A sky130_fd_sc_hd__inv_1_71/A
+ sky130_fd_sc_hd__nand2_8_3/Y sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_90 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_6 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_10/HI
+ sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_6/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# sky130_fd_sc_hd__dfbbn_1_6/a_557_413# sky130_fd_sc_hd__dfbbn_1_6/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_6/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__dfbbn_1_6/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_581_47# sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# sky130_fd_sc_hd__dfbbn_1_6/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# sky130_fd_sc_hd__dfbbn_1_6/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_4 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_4/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_48 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_37 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_39/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_26 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_27/Y
+ sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_15 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_15/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_59 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__inv_1_59/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_8_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__nand2_8_3/Y
+ sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_91 V_GND sky130_fd_sc_hd__fill_4_84/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 V_GND sky130_fd_sc_hd__fill_4_72/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_7 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF16.Q
+ sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_12/HI
+ sky130_fd_sc_hd__inv_1_17/Y FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# sky130_fd_sc_hd__dfbbn_1_7/a_557_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# sky130_fd_sc_hd__dfbbn_1_7/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_581_47# sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# sky130_fd_sc_hd__dfbbn_1_7/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# sky130_fd_sc_hd__dfbbn_1_7/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_5 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_5/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_49 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_38 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_40/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_27 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_28/Y
+ sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_16 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_16/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_8_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_64/A
+ sky130_fd_sc_hd__inv_1_93/A sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_92 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 V_GND sky130_fd_sc_hd__fill_4_73/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_70 V_GND sky130_fd_sc_hd__fill_4_69/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_8 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_13/HI
+ sky130_fd_sc_hd__inv_1_18/Y FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__dfbbn_1_8/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_8/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# sky130_fd_sc_hd__dfbbn_1_8/a_557_413# sky130_fd_sc_hd__dfbbn_1_8/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_8/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# sky130_fd_sc_hd__dfbbn_1_8/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_581_47# sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# sky130_fd_sc_hd__dfbbn_1_8/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# sky130_fd_sc_hd__dfbbn_1_8/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_6 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_6/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_39 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_39/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_28 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_33/Y
+ sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_17 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF16.Q
+ sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_8_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_68/A
+ sky130_fd_sc_hd__inv_1_70/A sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_60 V_GND sky130_fd_sc_hd__fill_4_63/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 V_GND sky130_fd_sc_hd__fill_4_68/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 V_GND sky130_fd_sc_hd__fill_4_74/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 V_GND sky130_fd_sc_hd__fill_4_87/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_9 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_11/HI
+ sky130_fd_sc_hd__inv_1_19/Y FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_9/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# sky130_fd_sc_hd__dfbbn_1_9/a_557_413# sky130_fd_sc_hd__dfbbn_1_9/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# sky130_fd_sc_hd__dfbbn_1_9/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_581_47# sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# sky130_fd_sc_hd__dfbbn_1_9/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# sky130_fd_sc_hd__dfbbn_1_9/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_7 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_7/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_29 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_32/Y
+ sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_18 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_8_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_93/A
+ sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_50 V_GND sky130_fd_sc_hd__fill_4_60/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 V_GND sky130_fd_sc_hd__fill_4_58/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_72 V_GND sky130_fd_sc_hd__fill_4_74/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 V_GND sky130_fd_sc_hd__fill_4_69/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 V_GND sky130_fd_sc_hd__fill_4_85/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_8 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_8/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_19 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__inv_1_19/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_8_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_70/A
+ sky130_fd_sc_hd__inv_1_68/A sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_95 V_GND sky130_fd_sc_hd__fill_4_87/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 V_GND sky130_fd_sc_hd__fill_4_63/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_62 V_GND sky130_fd_sc_hd__fill_4_56/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 V_GND sky130_fd_sc_hd__fill_4_72/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_73 V_GND sky130_fd_sc_hd__fill_4_73/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_40 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_9 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_9/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor2_1_0 V_GND V_LOW V_GND V_LOW Reset CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nor2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nand2_8_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand3_1_0/Y CLOCK_GEN.SR_Op.Q
+ sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_96 V_GND sky130_fd_sc_hd__fill_4_85/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_63 V_GND sky130_fd_sc_hd__fill_4_60/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_52 V_GND sky130_fd_sc_hd__fill_4_63/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 V_GND sky130_fd_sc_hd__fill_4_75/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 V_GND sky130_fd_sc_hd__fill_4_68/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_110 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_8_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_63/Y sky130_fd_sc_hd__nand2_8_9/Y
+ CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__decap_4_20 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_97 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_53 V_GND sky130_fd_sc_hd__fill_4_56/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 V_GND sky130_fd_sc_hd__fill_4_73/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 V_GND sky130_fd_sc_hd__fill_4_68/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_100 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__inv_1_100/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_111 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_54 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_10 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 V_GND sky130_fd_sc_hd__fill_4_56/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 V_GND sky130_fd_sc_hd__fill_4_73/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_76 V_GND sky130_fd_sc_hd__fill_4_68/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_50 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_51/HI
+ sky130_fd_sc_hd__inv_1_49/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_50/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_50/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# sky130_fd_sc_hd__dfbbn_1_50/a_557_413# sky130_fd_sc_hd__dfbbn_1_50/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_50/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# sky130_fd_sc_hd__dfbbn_1_50/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_581_47# sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# sky130_fd_sc_hd__dfbbn_1_50/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_50/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_101 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__inv_1_101/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_112 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__inv_1_112/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_99 V_GND sky130_fd_sc_hd__fill_4_84/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_11 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_88 V_GND sky130_fd_sc_hd__fill_4_75/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 V_GND sky130_fd_sc_hd__fill_4_72/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_77 V_GND sky130_fd_sc_hd__fill_4_69/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_160 V_GND sky130_fd_sc_hd__fill_8_819/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_40 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_47/HI
+ sky130_fd_sc_hd__inv_1_109/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_40/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_40/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# sky130_fd_sc_hd__dfbbn_1_40/a_557_413# sky130_fd_sc_hd__dfbbn_1_40/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_40/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# sky130_fd_sc_hd__dfbbn_1_40/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_581_47# sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# sky130_fd_sc_hd__dfbbn_1_40/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_40/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_51 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_40/HI
+ sky130_fd_sc_hd__inv_1_48/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_51/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__dfbbn_1_51/a_557_413# sky130_fd_sc_hd__dfbbn_1_51/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_51/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__dfbbn_1_51/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_581_47# sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# sky130_fd_sc_hd__dfbbn_1_51/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_51/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_102 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__inv_1_102/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_113 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_85/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_45 V_GND sky130_fd_sc_hd__fill_4_60/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_12 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_89 V_GND sky130_fd_sc_hd__fill_4_75/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 V_GND sky130_fd_sc_hd__fill_4_74/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_78 V_GND sky130_fd_sc_hd__fill_4_74/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_150 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_161 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_30 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_41/HI
+ sky130_fd_sc_hd__inv_1_102/Y FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__dfbbn_1_30/a_557_413# sky130_fd_sc_hd__dfbbn_1_30/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_581_47# sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# sky130_fd_sc_hd__dfbbn_1_30/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_41 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_27/HI
+ sky130_fd_sc_hd__inv_1_112/Y RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_41/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_41/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# sky130_fd_sc_hd__dfbbn_1_41/a_557_413# sky130_fd_sc_hd__dfbbn_1_41/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_41/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# sky130_fd_sc_hd__dfbbn_1_41/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_581_47# sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# sky130_fd_sc_hd__dfbbn_1_41/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_41/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_103 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__inv_1_103/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_114 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_1_72/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_13 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_46 V_GND sky130_fd_sc_hd__fill_4_63/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 V_GND sky130_fd_sc_hd__fill_4_56/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_79 V_GND sky130_fd_sc_hd__fill_4_75/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_68 V_GND sky130_fd_sc_hd__fill_4_69/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_140 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_151 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_31 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_35/HI
+ sky130_fd_sc_hd__inv_1_101/Y FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_31/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_31/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__dfbbn_1_31/a_557_413# sky130_fd_sc_hd__dfbbn_1_31/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_31/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__dfbbn_1_31/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_581_47# sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# sky130_fd_sc_hd__dfbbn_1_31/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_31/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_42 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_29/HI
+ sky130_fd_sc_hd__inv_1_59/Y RISING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_42/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__dfbbn_1_42/a_557_413# sky130_fd_sc_hd__dfbbn_1_42/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# sky130_fd_sc_hd__dfbbn_1_42/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_581_47# sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# sky130_fd_sc_hd__dfbbn_1_42/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_42/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_20 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_20/HI
+ sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__dfbbn_1_20/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_20/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# sky130_fd_sc_hd__dfbbn_1_20/a_557_413# sky130_fd_sc_hd__dfbbn_1_20/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__dfbbn_1_20/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# sky130_fd_sc_hd__dfbbn_1_20/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_581_47# sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# sky130_fd_sc_hd__dfbbn_1_20/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_20/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_104 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_115 V_GND V_HIGH V_GND V_HIGH Reset transmission_gate_0/GN
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_14 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_36 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 V_GND sky130_fd_sc_hd__fill_4_60/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 V_GND sky130_fd_sc_hd__fill_4_72/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_141 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_130 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_152 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_2_0 V_GND V_HIGH V_HIGH V_GND sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_2_0/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__dfbbn_1_32 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_39/HI
+ sky130_fd_sc_hd__inv_1_100/Y FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_32/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# sky130_fd_sc_hd__dfbbn_1_32/a_557_413# sky130_fd_sc_hd__dfbbn_1_32/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_32/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# sky130_fd_sc_hd__dfbbn_1_32/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_581_47# sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# sky130_fd_sc_hd__dfbbn_1_32/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_32/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_43 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_50/HI
+ sky130_fd_sc_hd__inv_1_90/Y RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__dfbbn_1_43/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# sky130_fd_sc_hd__dfbbn_1_43/a_557_413# sky130_fd_sc_hd__dfbbn_1_43/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# sky130_fd_sc_hd__dfbbn_1_43/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_581_47# sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# sky130_fd_sc_hd__dfbbn_1_43/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_21 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_26/HI
+ sky130_fd_sc_hd__inv_1_58/Y RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_21/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_21/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# sky130_fd_sc_hd__dfbbn_1_21/a_557_413# sky130_fd_sc_hd__dfbbn_1_21/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_21/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__dfbbn_1_21/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_581_47# sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# sky130_fd_sc_hd__dfbbn_1_21/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_21/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_10 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF18.Q
+ sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_14/HI
+ sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_10/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# sky130_fd_sc_hd__dfbbn_1_10/a_557_413# sky130_fd_sc_hd__dfbbn_1_10/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_10/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# sky130_fd_sc_hd__dfbbn_1_10/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_581_47# sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# sky130_fd_sc_hd__dfbbn_1_10/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_10/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_105 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__inv_1_105/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_116 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_48 V_GND sky130_fd_sc_hd__fill_4_58/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 V_GND sky130_fd_sc_hd__fill_4_58/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_15 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xtransmission_gate_0 Reset V_HIGH V_GND V_SENSE transmission_gate_0/GN transmission_gate
Xsky130_fd_sc_hd__decap_4_142 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_120 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_131 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_153 V_GND sky130_fd_sc_hd__fill_8_819/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_33 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_37/HI
+ sky130_fd_sc_hd__inv_1_98/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__dfbbn_1_33/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# sky130_fd_sc_hd__dfbbn_1_33/a_557_413# sky130_fd_sc_hd__dfbbn_1_33/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_581_47# sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# sky130_fd_sc_hd__dfbbn_1_33/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_22 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_32/HI
+ sky130_fd_sc_hd__inv_1_61/Y RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__dfbbn_1_22/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_22/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# sky130_fd_sc_hd__dfbbn_1_22/a_557_413# sky130_fd_sc_hd__dfbbn_1_22/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_22/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__dfbbn_1_22/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_581_47# sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# sky130_fd_sc_hd__dfbbn_1_22/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_22/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_11 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF17.Q
+ sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_16/HI
+ sky130_fd_sc_hd__inv_1_23/Y FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__dfbbn_1_11/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_11/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_581_47# sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# sky130_fd_sc_hd__dfbbn_1_11/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_11/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_44 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_24/HI
+ sky130_fd_sc_hd__inv_1_111/Y RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_44/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# sky130_fd_sc_hd__dfbbn_1_44/a_557_413# sky130_fd_sc_hd__dfbbn_1_44/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# sky130_fd_sc_hd__dfbbn_1_44/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_581_47# sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# sky130_fd_sc_hd__dfbbn_1_44/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_106 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__inv_1_106/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_117 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__inv_1_119/Y
+ sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__conb_1_50 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_50/LO
+ sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_16 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 V_GND sky130_fd_sc_hd__fill_4_58/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_38 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_110 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_143 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_132 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_121 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_154 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_34 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_44/HI
+ sky130_fd_sc_hd__inv_1_110/Y FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__dfbbn_1_34/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_34/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__dfbbn_1_34/a_557_413# sky130_fd_sc_hd__dfbbn_1_34/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_34/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# sky130_fd_sc_hd__dfbbn_1_34/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# sky130_fd_sc_hd__dfbbn_1_34/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_34/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_45 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_48/HI
+ sky130_fd_sc_hd__inv_1_108/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_45/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# sky130_fd_sc_hd__dfbbn_1_45/a_557_413# sky130_fd_sc_hd__dfbbn_1_45/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# sky130_fd_sc_hd__dfbbn_1_45/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_581_47# sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# sky130_fd_sc_hd__dfbbn_1_45/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__dfbbn_1_45/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_23 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_31/HI
+ sky130_fd_sc_hd__inv_1_62/Y RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# sky130_fd_sc_hd__dfbbn_1_23/a_557_413# sky130_fd_sc_hd__dfbbn_1_23/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# sky130_fd_sc_hd__dfbbn_1_23/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_12 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF19.Q
+ sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_17/HI
+ sky130_fd_sc_hd__inv_1_22/Y FULL_COUNTER.COUNT_SUB_DFF18.Q sky130_fd_sc_hd__dfbbn_1_12/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# sky130_fd_sc_hd__dfbbn_1_12/a_557_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_581_47# sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# sky130_fd_sc_hd__dfbbn_1_12/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_107 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__inv_1_107/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_118 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__nand3_1_2/B
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__conb_1_40 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_40/LO
+ sky130_fd_sc_hd__conb_1_40/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_51 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_51/LO
+ sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_17 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_144 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_111 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_122 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_133 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_100 V_GND sky130_fd_sc_hd__fill_4_87/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_155 V_GND sky130_fd_sc_hd__fill_8_819/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_46 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_36/HI
+ sky130_fd_sc_hd__inv_1_99/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__dfbbn_1_46/a_557_413# sky130_fd_sc_hd__dfbbn_1_46/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_581_47# sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# sky130_fd_sc_hd__dfbbn_1_46/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_35 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_43/HI
+ sky130_fd_sc_hd__inv_1_105/Y FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_35/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# sky130_fd_sc_hd__dfbbn_1_35/a_557_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_581_47# sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# sky130_fd_sc_hd__dfbbn_1_35/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_24 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_28/HI
+ sky130_fd_sc_hd__inv_1_60/Y RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__dfbbn_1_24/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__dfbbn_1_24/a_557_413# sky130_fd_sc_hd__dfbbn_1_24/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__dfbbn_1_24/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_581_47# sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# sky130_fd_sc_hd__dfbbn_1_24/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_13 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_6/HI
+ sky130_fd_sc_hd__inv_1_12/Y FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__dfbbn_1_13/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__dfbbn_1_13/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# sky130_fd_sc_hd__dfbbn_1_13/a_557_413# sky130_fd_sc_hd__dfbbn_1_13/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__dfbbn_1_13/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_581_47# sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# sky130_fd_sc_hd__dfbbn_1_13/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_108 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__inv_1_108/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_119 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_119/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__conb_1_41 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_41/LO
+ sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_30 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_30/LO
+ sky130_fd_sc_hd__conb_1_30/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand3_1_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_66/Y
+ sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__nand3_1_0/a_193_47#
+ sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_18 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_29 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_112 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_101 V_GND sky130_fd_sc_hd__fill_4_84/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_123 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_145 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_134 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_156 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_36 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_42/HI
+ sky130_fd_sc_hd__inv_1_104/Y FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_36/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__dfbbn_1_36/a_557_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# sky130_fd_sc_hd__dfbbn_1_36/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_25 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_22/HI
+ sky130_fd_sc_hd__inv_1_53/Y RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_25/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# sky130_fd_sc_hd__dfbbn_1_25/a_557_413# sky130_fd_sc_hd__dfbbn_1_25/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_581_47# sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# sky130_fd_sc_hd__dfbbn_1_25/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_47 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_25/HI
+ sky130_fd_sc_hd__inv_1_57/Y RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_47/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# sky130_fd_sc_hd__dfbbn_1_47/a_557_413# sky130_fd_sc_hd__dfbbn_1_47/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# sky130_fd_sc_hd__dfbbn_1_47/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_581_47# sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__dfbbn_1_47/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_14 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_18/HI
+ sky130_fd_sc_hd__inv_1_15/Y FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_14/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__dfbbn_1_14/a_557_413# sky130_fd_sc_hd__dfbbn_1_14/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_581_47# sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# sky130_fd_sc_hd__dfbbn_1_14/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_109 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__conb_1_42 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_42/LO
+ sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_31 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_31/LO
+ sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_20 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_20/LO
+ sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand3_1_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_94/Y
+ sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__nand3_1_1/a_193_47#
+ sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_19 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_146 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_113 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_102 V_GND sky130_fd_sc_hd__fill_4_85/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_124 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_135 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_157 V_GND sky130_fd_sc_hd__fill_8_819/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_15 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_15/HI
+ sky130_fd_sc_hd__inv_1_20/Y FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# sky130_fd_sc_hd__dfbbn_1_15/a_557_413# sky130_fd_sc_hd__dfbbn_1_15/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__dfbbn_1_15/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_581_47# sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# sky130_fd_sc_hd__dfbbn_1_15/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_37 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_45/HI
+ sky130_fd_sc_hd__inv_1_103/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__dfbbn_1_37/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# sky130_fd_sc_hd__dfbbn_1_37/a_557_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_581_47# sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# sky130_fd_sc_hd__dfbbn_1_37/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_48 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__dfbbn_1_48/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_34/HI
+ sky130_fd_sc_hd__inv_1_88/Y RISING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_48/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# sky130_fd_sc_hd__dfbbn_1_48/a_557_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_381_47# sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_581_47# sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# sky130_fd_sc_hd__dfbbn_1_48/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_26 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_30/HI
+ sky130_fd_sc_hd__inv_1_55/Y RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__dfbbn_1_26/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# sky130_fd_sc_hd__dfbbn_1_26/a_557_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_581_47# sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# sky130_fd_sc_hd__dfbbn_1_26/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_43 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_43/LO
+ sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_32 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_32/LO
+ sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_21 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_21/LO
+ sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_10 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_10/LO
+ sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand3_1_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__nand3_1_2/B
+ sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand3_1_2/a_193_47#
+ sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_147 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_114 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_103 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_125 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_136 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_158 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_38 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_49/HI
+ sky130_fd_sc_hd__inv_1_106/Y FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__dfbbn_1_38/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_38/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# sky130_fd_sc_hd__dfbbn_1_38/a_557_413# sky130_fd_sc_hd__dfbbn_1_38/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_38/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# sky130_fd_sc_hd__dfbbn_1_38/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_581_47# sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# sky130_fd_sc_hd__dfbbn_1_38/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__dfbbn_1_38/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_49 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_38/HI
+ sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__dfbbn_1_49/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# sky130_fd_sc_hd__dfbbn_1_49/a_557_413# sky130_fd_sc_hd__dfbbn_1_49/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_581_47# sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# sky130_fd_sc_hd__dfbbn_1_49/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_27 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_23/HI
+ sky130_fd_sc_hd__inv_1_56/Y RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__dfbbn_1_27/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__dfbbn_1_27/a_557_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_581_47# sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# sky130_fd_sc_hd__dfbbn_1_27/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_16 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_4/HI
+ sky130_fd_sc_hd__inv_1_8/Y FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_16/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_16/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# sky130_fd_sc_hd__dfbbn_1_16/a_557_413# sky130_fd_sc_hd__dfbbn_1_16/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_16/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_581_47# sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# sky130_fd_sc_hd__dfbbn_1_16/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_22 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_22/LO
+ sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_11 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_11/LO
+ sky130_fd_sc_hd__conb_1_11/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_44 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_44/LO
+ sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_33 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_33/LO
+ sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_115 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_148 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_126 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_137 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_104 V_GND sky130_fd_sc_hd__fill_4_87/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_159 V_GND V_HIGH V_GND V_HIGH sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_39 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__dfbbn_1_39/Q_N sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_46/HI
+ sky130_fd_sc_hd__inv_1_107/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__dfbbn_1_39/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_791_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# sky130_fd_sc_hd__dfbbn_1_39/a_557_413# sky130_fd_sc_hd__dfbbn_1_39/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_381_47# sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_581_47# sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# sky130_fd_sc_hd__dfbbn_1_39/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_28 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_21/HI
+ sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# sky130_fd_sc_hd__dfbbn_1_28/a_557_413# sky130_fd_sc_hd__dfbbn_1_28/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_581_47# sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# sky130_fd_sc_hd__dfbbn_1_28/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_17 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_19/HI
+ sky130_fd_sc_hd__inv_1_4/Y FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__dfbbn_1_17/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# sky130_fd_sc_hd__dfbbn_1_17/a_557_413# sky130_fd_sc_hd__dfbbn_1_17/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_581_47# sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# sky130_fd_sc_hd__dfbbn_1_17/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_45 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_45/LO
+ sky130_fd_sc_hd__conb_1_45/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_34 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_34/LO
+ sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_23 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_23/LO
+ sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_12 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_12/LO
+ sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_105 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_149 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_116 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_127 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_138 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_29 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_33/HI
+ sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__dfbbn_1_29/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_791_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# sky130_fd_sc_hd__dfbbn_1_29/a_557_413# sky130_fd_sc_hd__dfbbn_1_29/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__dfbbn_1_29/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__dfbbn_1_29/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_581_47# sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# sky130_fd_sc_hd__dfbbn_1_29/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__dfbbn_1_29/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__dfbbn_1_18 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_9/HI
+ sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# sky130_fd_sc_hd__dfbbn_1_18/a_557_413# sky130_fd_sc_hd__dfbbn_1_18/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_581_47# sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# sky130_fd_sc_hd__dfbbn_1_18/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_35 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_35/LO
+ sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_46 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_46/LO
+ sky130_fd_sc_hd__conb_1_46/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_24 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_24/LO
+ sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_13 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_13/LO
+ sky130_fd_sc_hd__conb_1_13/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_117 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_128 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_106 V_GND sky130_fd_sc_hd__fill_4_85/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_139 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfbbn_1_19 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF4.Q
+ sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_5/HI
+ sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_19/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# sky130_fd_sc_hd__dfbbn_1_19/a_557_413# sky130_fd_sc_hd__dfbbn_1_19/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_581_47# sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# sky130_fd_sc_hd__dfbbn_1_19/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_1672_329#
+ sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__conb_1_47 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_47/LO
+ sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_36 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_36/LO
+ sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_25 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_25/LO
+ sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_14 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_14/LO
+ sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_118 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_129 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_107 V_GND sky130_fd_sc_hd__fill_4_84/VPB V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_48 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_48/LO
+ sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_37 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_37/LO
+ sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_26 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_26/LO
+ sky130_fd_sc_hd__conb_1_26/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_15 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_15/LO
+ sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_119 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_108 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_90 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__inv_1_90/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__conb_1_38 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_38/LO
+ sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_27 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_27/LO
+ sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_16 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_16/LO
+ sky130_fd_sc_hd__conb_1_16/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_49 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_49/LO
+ sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_4_109 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_91 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_91/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_80 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__inv_1_96/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_39 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_39/LO
+ sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_28 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_28/LO
+ sky130_fd_sc_hd__conb_1_28/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_17 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_17/LO
+ sky130_fd_sc_hd__conb_1_17/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_1_92 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_97/Y sky130_fd_sc_hd__inv_1_92/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_81 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_81/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_70 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_70/A sky130_fd_sc_hd__inv_1_70/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_1/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_29 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_29/LO
+ sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_18 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_18/LO
+ sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__inv_1_82 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_91/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_60 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF8.Q
+ sky130_fd_sc_hd__inv_1_60/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_93 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_93/A sky130_fd_sc_hd__inv_1_93/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_71 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_71/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_2/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_19 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_19/LO
+ sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_1_0/Y
+ sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_50 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_50/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_83 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_86/Y sky130_fd_sc_hd__inv_1_83/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_61 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_94 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_94/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_72 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__inv_1_72/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__conb_1_3/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__nand2_1_2/A
+ sky130_fd_sc_hd__inv_1_75/A sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_84 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_89/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_51 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_51/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_62 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF9.Q
+ sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_73 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_75/A sky130_fd_sc_hd__inv_1_95/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_40 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_40/A sky130_fd_sc_hd__inv_1_44/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_95 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_95/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__conb_1_4/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_2/A
+ sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_85 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_85/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_74 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__inv_1_74/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_41 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_46/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_96 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_96/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_52 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF14.Q
+ sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_63 V_GND V_LOW V_GND V_LOW Reset sky130_fd_sc_hd__inv_1_63/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_30 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_31/Y
+ sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_5/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_3 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__nand2_1_3/Y
+ sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfbbn_1_0 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_1/HI
+ sky130_fd_sc_hd__inv_1_5/Y FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_0/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_0/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# sky130_fd_sc_hd__dfbbn_1_0/a_557_413# sky130_fd_sc_hd__dfbbn_1_0/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_0/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__dfbbn_1_0/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_581_47# sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# sky130_fd_sc_hd__dfbbn_1_0/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# sky130_fd_sc_hd__dfbbn_1_0/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_86 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_86/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_97 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__inv_1_97/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_75 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_75/A sky130_fd_sc_hd__inv_1_75/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_42 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_42/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_64 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_64/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_53 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF15.Q
+ sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_31 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_31/A
+ sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_20 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__inv_1_20/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_6 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_6/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_4 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__nand2_8_3/A
+ sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfbbn_1_1 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_2/HI
+ sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_1/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__dfbbn_1_1/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# sky130_fd_sc_hd__dfbbn_1_1/a_557_413# sky130_fd_sc_hd__dfbbn_1_1/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_1/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# sky130_fd_sc_hd__dfbbn_1_1/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_581_47# sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# sky130_fd_sc_hd__dfbbn_1_1/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# sky130_fd_sc_hd__dfbbn_1_1/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_32 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_32/A
+ sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_10 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_10/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_21 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF18.Q
+ sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_98 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF6.Q
+ sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_87 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_97/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_43 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_43/A sky130_fd_sc_hd__inv_1_43/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_76 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_94/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_65 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_54 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF13.Q
+ sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_7 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_7/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_1_5 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__nand2_1_5/Y
+ sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__dfbbn_1_2 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_3/HI
+ sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_119/Y sky130_fd_sc_hd__dfbbn_1_2/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_791_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_2/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# sky130_fd_sc_hd__dfbbn_1_2/a_557_413# sky130_fd_sc_hd__dfbbn_1_2/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__dfbbn_1_2/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# sky130_fd_sc_hd__dfbbn_1_2/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_581_47# sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# sky130_fd_sc_hd__dfbbn_1_2/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__dfbbn_1_2/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_0 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_44 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_45/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_55 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_66 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_66/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_33 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_2_0/Y
+ sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_11 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_22 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF19.Q
+ sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_99 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF7.Q
+ sky130_fd_sc_hd__inv_1_99/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_77 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_78/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_88 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF5.Q
+ sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_0/Y Reset
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_4_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_8 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__conb_1_8/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__dfbbn_1_3 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF1.Q
+ sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_0/HI
+ sky130_fd_sc_hd__inv_1_10/Y FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_791_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__dfbbn_1_3/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_581_47# sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__dfbbn_1_3/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__dfbbn_1_3/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_1 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_1/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_89 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_89/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_78 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_78/A sky130_fd_sc_hd__inv_1_79/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_45 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_45/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_56 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__inv_1_56/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_67 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_67/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_34 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_34/A
+ sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_12 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF10.Q
+ sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_23 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF17.Q
+ sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_1/Y Reset
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__decap_4_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_9 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__conb_1_9/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__nand2_8_0 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__nand3_1_2/B sky130_fd_sc_hd__inv_1_51/A
+ sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__dfbbn_1_4 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF11.Q
+ sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_7/HI
+ sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__dfbbn_1_4/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_4/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# sky130_fd_sc_hd__dfbbn_1_4/a_557_413# sky130_fd_sc_hd__dfbbn_1_4/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__dfbbn_1_4/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# sky130_fd_sc_hd__dfbbn_1_4/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_581_47# sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# sky130_fd_sc_hd__dfbbn_1_4/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# sky130_fd_sc_hd__dfbbn_1_4/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_2 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_79 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_80/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_35 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_75/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_46 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_46/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_57 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF2.Q
+ sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_68 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_68/A sky130_fd_sc_hd__inv_1_68/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_24 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_1/Y
+ sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_13 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_16_2 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_16_2/Y Reset
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__nand2_8_1 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_50/A
+ sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__nand2_8
Xsky130_fd_sc_hd__dfbbn_1_5 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF12.Q
+ sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_8/HI
+ sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__dfbbn_1_5/a_2136_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_891_329#
+ sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# sky130_fd_sc_hd__dfbbn_1_5/a_557_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21#
+ sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_581_47# sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# sky130_fd_sc_hd__dfbbn_1_5/a_1159_47#
+ sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# sky130_fd_sc_hd__dfbbn_1_5/a_27_47#
+ sky130_fd_sc_hd__dfbbn_1
Xsky130_fd_sc_hd__inv_1_3 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_14 V_GND V_LOW V_GND V_LOW FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_14/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_47 V_GND V_LOW V_GND V_LOW FALLING_COUNTER.COUNT_SUB_DFF0.Q
+ sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_36 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_43/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_58 V_GND V_LOW V_GND V_LOW RISING_COUNTER.COUNT_SUB_DFF3.Q
+ sky130_fd_sc_hd__inv_1_58/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_69 V_GND V_LOW V_GND V_LOW sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__inv_1_69/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_25 V_GND V_SENSE V_GND V_SENSE sky130_fd_sc_hd__inv_1_26/Y
+ sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1
C0 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__inv_1_57/Y 8.71e-19
C1 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__inv_1_22/Y 1.93e-21
C2 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__inv_16_1/Y 0.0018f
C3 sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__inv_1_60/Y 0.00158f
C4 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_70/A 0.045f
C5 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 3.05e-19
C6 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__inv_16_2/Y 0.00121f
C7 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0.00106f
C8 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 7.96e-20
C9 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 2.71e-19
C10 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__inv_1_102/Y 1.49e-20
C11 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 0.00207f
C12 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# V_LOW 0.0026f
C13 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/Q_N 1.89e-19
C14 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00114f
C15 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# V_LOW 0.00449f
C16 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00161f
C17 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_4/HI 0.0195f
C18 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 5.74e-19
C19 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 3.13e-21
C20 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 9.65e-21
C21 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 0.0036f
C22 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 5.82e-20
C23 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_1_5/Y 0.0064f
C24 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# V_GND 1.92e-19
C25 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# 0.00228f
C26 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 5.97e-20
C27 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 4.97e-19
C28 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# 8.67e-19
C29 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_105/Y 2.17e-21
C30 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0338f
C31 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# sky130_fd_sc_hd__inv_1_107/Y 0.00235f
C32 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_2/HI 0.103f
C33 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.49e-19
C34 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 0.0784f
C35 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__conb_1_31/HI 0.00225f
C36 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# V_GND -0.00441f
C37 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_72/A 0.0233f
C38 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__conb_1_0/HI 8.47e-19
C39 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__conb_1_1/HI 0.0144f
C40 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# V_GND 4.15e-19
C41 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.92e-20
C42 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_36/HI 0.0222f
C43 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__inv_1_103/Y 0.00596f
C44 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# -3.46e-20
C45 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__conb_1_19/HI 1.16e-20
C46 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_50/Y 7.63e-19
C47 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 8.66e-19
C48 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 1.18f
C49 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.49e-19
C50 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# sky130_fd_sc_hd__inv_1_61/Y 7.97e-21
C51 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 0.0235f
C52 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_30/HI 2.22e-19
C53 sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# sky130_fd_sc_hd__conb_1_34/HI 4.53e-19
C54 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_66/Y 1.08e-19
C55 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00283f
C56 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__conb_1_42/HI 0.00294f
C57 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__conb_1_45/HI 4.86e-20
C58 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__conb_1_5/LO 0.00187f
C59 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.5e-20
C60 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 0.00117f
C61 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__inv_1_59/Y 2.6e-20
C62 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__conb_1_24/HI -0.00776f
C63 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.067f
C64 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0.0326f
C65 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 6.39e-19
C66 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00297f
C67 sky130_fd_sc_hd__inv_1_64/A V_GND 0.146f
C68 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# -9.32e-20
C69 Reset RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0215f
C70 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_65/Y 3.53e-19
C71 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.104f
C72 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.6e-20
C73 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# -2.01e-20
C74 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# -0.00222f
C75 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.34e-22
C76 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_1_102/Y 3.91e-19
C77 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/Q_N -9.56e-20
C78 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 1.52e-19
C79 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 5.48e-21
C80 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_56/Y 0.00742f
C81 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -3.86e-20
C82 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 5.36e-22
C83 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_1_108/Y 0.00171f
C84 sky130_fd_sc_hd__dfbbn_1_15/Q_N FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00373f
C85 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 3.54e-21
C86 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__inv_1_4/Y 0.0107f
C87 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 1.28e-20
C88 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 9.61e-19
C89 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 1.15e-20
C90 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# V_LOW 0.00133f
C91 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_20/Y 7.45e-20
C92 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 5.9e-21
C93 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 8.06e-20
C94 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 2.61e-19
C95 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00107f
C96 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.52e-20
C97 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/Q_N 7.75e-19
C98 sky130_fd_sc_hd__inv_1_66/Y V_GND 0.118f
C99 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__nand2_8_9/Y 0.0196f
C100 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__nand3_1_2/B 1.4e-21
C101 sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__inv_1_75/A 1.7e-19
C102 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_57/Y 0.104f
C103 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 4.36e-19
C104 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.52e-19
C105 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# sky130_fd_sc_hd__conb_1_5/HI 0.00107f
C106 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 6.86e-20
C107 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 4.04e-21
C108 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 4.04e-21
C109 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_37/HI 3.73e-19
C110 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_45/A 0.0133f
C111 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# V_LOW -6.55e-19
C112 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 5.31e-19
C113 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 1.1e-20
C114 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 8.43e-20
C115 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# sky130_fd_sc_hd__conb_1_4/HI 1.47e-19
C116 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__conb_1_42/HI 3.27e-19
C117 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_103/Y 0.00463f
C118 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.571f
C119 sky130_fd_sc_hd__inv_1_106/Y V_GND 0.0699f
C120 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_16_2/Y 0.00335f
C121 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_95/Y 1.11e-19
C122 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# V_LOW 0.0272f
C123 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_102/Y 3.43e-20
C124 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__conb_1_37/LO 5.27e-20
C125 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 0.123f
C126 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# sky130_fd_sc_hd__inv_1_107/Y 2.12e-19
C127 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_67/Y 0.325f
C128 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0514f
C129 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 0.0214f
C130 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_10/HI 9.34e-20
C131 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.15e-19
C132 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# V_LOW -8.36e-19
C133 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_10/HI 5.23e-19
C134 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__conb_1_31/HI 0.00213f
C135 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# V_GND -0.00163f
C136 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__conb_1_9/HI -0.00392f
C137 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# -0.00263f
C138 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# -5.54e-21
C139 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__conb_1_10/HI 4.24e-19
C140 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__conb_1_36/HI -4.53e-19
C141 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__conb_1_36/HI 7.99e-19
C142 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_74/Y 7.42e-21
C143 sky130_fd_sc_hd__inv_1_12/Y V_GND 0.139f
C144 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__nand3_1_1/Y 0.0141f
C145 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_22/Y 0.00139f
C146 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.09e-20
C147 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_473_413# 2.14e-19
C148 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 1.81e-19
C149 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nor2_1_0/Y 0.0437f
C150 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0393f
C151 sky130_fd_sc_hd__inv_1_17/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0228f
C152 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__conb_1_11/HI -0.0122f
C153 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__inv_1_55/Y 1.28e-20
C154 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# V_LOW 0.00918f
C155 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# V_GND 0.00647f
C156 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# V_LOW 0.0234f
C157 sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# sky130_fd_sc_hd__conb_1_45/HI 0.00196f
C158 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.332f
C159 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.47e-19
C160 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__conb_1_32/HI 2.25e-20
C161 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__inv_1_59/Y 1.55e-19
C162 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__inv_1_10/Y 0.00459f
C163 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# V_GND -0.0071f
C164 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__conb_1_13/HI 7.93e-19
C165 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# sky130_fd_sc_hd__conb_1_24/HI 2.62e-20
C166 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__conb_1_40/HI 2.81e-20
C167 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 0.0402f
C168 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 5.4e-19
C169 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 1.59e-22
C170 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 5.45e-19
C171 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/Q_N -4.33e-20
C172 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 1.92e-21
C173 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nor2_1_0/Y 3.05e-19
C174 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_23/Y 0.00316f
C175 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__nand3_1_1/Y 0.0073f
C176 Reset sky130_fd_sc_hd__inv_1_76/A 0.0272f
C177 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# -9.32e-20
C178 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0209f
C179 sky130_fd_sc_hd__fill_4_75/VPB V_LOW 0.797f
C180 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 7.43e-19
C181 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.00839f
C182 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF3.Q 0.11f
C183 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 8.26e-21
C184 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.62e-20
C185 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00965f
C186 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# V_GND 0.0059f
C187 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# V_GND 0.00525f
C188 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__nand2_1_0/Y 0.00132f
C189 sky130_fd_sc_hd__nand3_1_1/Y V_GND 0.208f
C190 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 7.62e-19
C191 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# V_GND -0.0463f
C192 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_112/Y 1.16e-19
C193 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# sky130_fd_sc_hd__inv_1_21/Y 2.63e-19
C194 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.375f
C195 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 5.96e-19
C196 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 0.00226f
C197 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# V_LOW 9.26e-19
C198 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_107/Y 6.11e-20
C199 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 2.5e-19
C200 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_12/HI 7.11e-19
C201 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -5.54e-21
C202 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# -2.14e-19
C203 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# 6.85e-20
C204 sky130_fd_sc_hd__dfbbn_1_38/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.12e-21
C205 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_16_1/Y 4.85e-21
C206 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 8.14e-21
C207 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_62/Y 1.01e-19
C208 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0.00114f
C209 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 0.0116f
C210 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 4.03e-19
C211 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.00278f
C212 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 0.0116f
C213 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__conb_1_22/HI 3.71e-19
C214 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_76/A 1.84e-19
C215 sky130_fd_sc_hd__dfbbn_1_32/Q_N V_LOW -0.00461f
C216 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_46/HI 4.56e-21
C217 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0786f
C218 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# 6.68e-21
C219 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# sky130_fd_sc_hd__conb_1_42/HI -0.00236f
C220 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 9.19e-22
C221 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 1.38e-20
C222 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__inv_1_90/Y 1.2e-19
C223 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 1.16e-19
C224 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# V_GND -0.00433f
C225 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_891_329# -0.00159f
C226 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# -0.00882f
C227 sky130_fd_sc_hd__inv_1_2/A V_GND 0.0167f
C228 sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# V_LOW 2.94e-20
C229 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.88e-19
C230 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# V_LOW 0.00955f
C231 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_5/HI 0.00134f
C232 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# 0.0456f
C233 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.00261f
C234 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 0.00115f
C235 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.08e-21
C236 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# V_LOW -0.00389f
C237 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_50/Y 0.00135f
C238 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.35e-19
C239 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# -9.32e-20
C240 sky130_fd_sc_hd__inv_1_47/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0914f
C241 Reset sky130_fd_sc_hd__inv_1_112/Y 0.00463f
C242 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_58/Y 2.47e-19
C243 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# sky130_fd_sc_hd__conb_1_36/HI -0.00109f
C244 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.101f
C245 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# V_LOW 0.00318f
C246 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_19/LO 0.0486f
C247 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# 1.19e-20
C248 sky130_fd_sc_hd__nand2_1_5/a_113_47# sky130_fd_sc_hd__inv_1_80/A 6.28e-21
C249 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 2.86e-20
C250 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00159f
C251 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.00194f
C252 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__inv_16_0/Y 0.0212f
C253 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 1.97e-22
C254 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# V_GND 7.24e-19
C255 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# V_LOW -0.00266f
C256 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# V_GND 2.59e-19
C257 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# -0.00482f
C258 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_891_329# -2.2e-20
C259 sky130_fd_sc_hd__inv_1_47/Y V_LOW 0.0633f
C260 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1_0/Y 5.73e-19
C261 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# -6.43e-19
C262 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# -0.0185f
C263 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 7e-19
C264 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# V_GND 7.04e-19
C265 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 3.2e-21
C266 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 5.3e-21
C267 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__inv_1_10/Y 1.07e-21
C268 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# V_GND -0.00992f
C269 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__conb_1_13/HI -0.00426f
C270 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 5.49e-20
C271 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# V_LOW 9.11e-19
C272 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00331f
C273 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_45/Y 6.18e-21
C274 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__conb_1_24/HI 7.43e-21
C275 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_381_47# -0.00144f
C276 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__conb_1_40/HI 9.37e-20
C277 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/Q_N 0.0249f
C278 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# -0.00519f
C279 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# V_GND 0.00212f
C280 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# V_GND -0.172f
C281 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/Q_N -4.33e-20
C282 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 8.72e-22
C283 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.13e-20
C284 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_80/A 0.236f
C285 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 6.19e-20
C286 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0.00611f
C287 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0.00622f
C288 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0251f
C289 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_381_47# 1.9e-19
C290 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# Reset 5.39e-19
C291 sky130_fd_sc_hd__conb_1_49/LO sky130_fd_sc_hd__inv_16_1/Y 0.0929f
C292 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0131f
C293 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# V_GND -6.34e-19
C294 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_68/A 3.27e-19
C295 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# V_GND 4.66e-19
C296 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# V_LOW 0.00652f
C297 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__conb_1_44/HI 0.00158f
C298 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF9.Q 9.04e-19
C299 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_83/Y 4.49e-19
C300 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_56/Y 1.43e-19
C301 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_193_47# 0.0297f
C302 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# V_LOW 1.38e-19
C303 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# V_GND 3.78e-19
C304 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__conb_1_36/LO 0.0121f
C305 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# V_LOW -0.00389f
C306 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_51/HI 0.177f
C307 sky130_fd_sc_hd__nand2_8_3/Y V_GND -0.00576f
C308 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF2.Q 9.11e-20
C309 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.009f
C310 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.89e-19
C311 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_40/A 4.26e-19
C312 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# 2.86e-19
C313 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 6.34e-19
C314 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 7.88e-21
C315 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# V_GND 5.15e-19
C316 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_13/Y 0.00314f
C317 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 4.8e-19
C318 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# sky130_fd_sc_hd__inv_16_1/Y 3.08e-20
C319 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 1.24e-19
C320 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__inv_1_101/Y 2.2e-19
C321 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# -9.32e-20
C322 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 9.25e-20
C323 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# -8.01e-19
C324 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_941_21# -0.0116f
C325 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# Reset 0.00135f
C326 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 5.71e-21
C327 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# V_GND 3.67e-19
C328 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_557_413# 0.0023f
C329 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__inv_1_21/Y 3.09e-21
C330 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# V_GND 0.00103f
C331 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 8.85e-19
C332 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_557_413# -0.0012f
C333 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# -0.00335f
C334 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# V_GND 6.73e-19
C335 FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_46/HI 0.0697f
C336 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0396f
C337 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__inv_1_90/Y 1.33e-19
C338 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# V_LOW -0.00261f
C339 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.62e-19
C340 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# V_GND 0.00529f
C341 FALLING_COUNTER.COUNT_SUB_DFF4.Q Reset 0.886f
C342 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# -0.00385f
C343 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 1.26e-20
C344 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 2.89e-20
C345 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 2.89e-20
C346 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0148f
C347 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__conb_1_2/HI 1.57e-19
C348 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.44e-19
C349 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# V_LOW 0.00185f
C350 sky130_fd_sc_hd__conb_1_24/LO V_GND 0.00261f
C351 sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF15.Q 6.71e-21
C352 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.21e-21
C353 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# -0.00887f
C354 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_891_329# -0.00161f
C355 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.027f
C356 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/Q_N -4.24e-20
C357 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__conb_1_44/HI 0.0152f
C358 sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__inv_2_0/Y 0.0146f
C359 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__conb_1_47/HI 0.00101f
C360 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# V_LOW 3.56e-20
C361 sky130_fd_sc_hd__conb_1_46/LO V_GND -3.53e-19
C362 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_381_47# 9.87e-20
C363 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# V_GND 2.94e-19
C364 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 1.59e-19
C365 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.16e-19
C366 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__inv_1_5/Y 5.2e-20
C367 RISING_COUNTER.COUNT_SUB_DFF12.Q V_GND 4.39f
C368 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0335f
C369 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.25e-19
C370 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# sky130_fd_sc_hd__inv_1_12/Y 2.28e-19
C371 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__inv_1_65/Y 7.25e-19
C372 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 1.67e-19
C373 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 1.6e-20
C374 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# sky130_fd_sc_hd__inv_1_12/Y 0.00106f
C375 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# -0.00142f
C376 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0155f
C377 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 8.64e-19
C378 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_16/LO 8.84e-20
C379 sky130_fd_sc_hd__conb_1_46/LO sky130_fd_sc_hd__inv_1_106/Y 0.122f
C380 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# -6.8e-19
C381 FULL_COUNTER.COUNT_SUB_DFF9.Q V_LOW 3.33f
C382 sky130_fd_sc_hd__conb_1_35/LO V_GND -0.00433f
C383 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_791_47# 1.64e-21
C384 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# sky130_fd_sc_hd__inv_1_9/Y 3.02e-21
C385 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0.00343f
C386 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# V_LOW 0.0125f
C387 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.84e-19
C388 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# -1.44e-20
C389 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.88e-19
C390 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# V_LOW 4.61e-20
C391 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_74/Y 6.68e-19
C392 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_581_47# -7.91e-19
C393 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_68/A 0.0809f
C394 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_70/A 1.75e-20
C395 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 2.74e-19
C396 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 0.00174f
C397 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# V_GND -0.00108f
C398 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# V_LOW 0.00592f
C399 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# V_GND 1.97e-19
C400 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 2.44e-20
C401 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# 2.55e-22
C402 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# 2.61e-21
C403 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.84e-20
C404 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 0.00893f
C405 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.041f
C406 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0143f
C407 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# -2.65e-20
C408 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 7.95e-19
C409 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 6.37e-20
C410 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 2.44e-19
C411 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -6.23e-21
C412 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_381_47# -0.00472f
C413 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_78/A 0.00355f
C414 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__conb_1_36/LO 9.67e-19
C415 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.98e-21
C416 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_791_47# -6.51e-19
C417 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 8.87e-20
C418 sky130_fd_sc_hd__inv_1_53/Y V_LOW 0.312f
C419 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0865f
C420 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# V_GND 0.0244f
C421 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__conb_1_36/LO 4.7e-20
C422 sky130_fd_sc_hd__nand2_8_4/a_27_47# V_LOW -0.00661f
C423 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.8e-20
C424 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# V_GND -0.00527f
C425 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_6/HI 0.0116f
C426 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_5/Y 0.00206f
C427 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.57e-20
C428 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_75/A 6.28e-21
C429 sky130_fd_sc_hd__conb_1_2/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 0.258f
C430 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 2.43e-21
C431 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__inv_1_13/Y 1.22e-21
C432 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 6.07e-20
C433 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00466f
C434 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# V_GND 3.29e-19
C435 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__conb_1_47/LO 1.29e-19
C436 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__inv_1_20/Y 7.56e-20
C437 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/Q_N -4.78e-20
C438 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_97/A 1.8e-19
C439 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 6.17e-19
C440 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_647_21# -0.00631f
C441 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_473_413# -3.06e-20
C442 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# -1.76e-19
C443 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# -7.17e-20
C444 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_18/LO 0.00496f
C445 sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__inv_1_100/Y 0.0594f
C446 sky130_fd_sc_hd__inv_1_110/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.87e-20
C447 sky130_fd_sc_hd__conb_1_14/LO FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00585f
C448 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 2.52e-19
C449 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 9.75e-19
C450 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 1.68e-19
C451 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 5.17e-21
C452 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.21e-19
C453 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0217f
C454 sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__conb_1_22/HI 0.00101f
C455 sky130_fd_sc_hd__conb_1_9/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 2.89e-20
C456 sky130_fd_sc_hd__conb_1_1/HI V_LOW 0.0379f
C457 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__conb_1_8/HI 5.66e-20
C458 sky130_fd_sc_hd__inv_1_88/Y Reset 0.0035f
C459 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_98/Y 1.84e-19
C460 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# Reset 5.13e-21
C461 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# -6.23e-21
C462 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# -3.04e-19
C463 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_1_6/Y 0.00728f
C464 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 0.026f
C465 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0047f
C466 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 4.28e-19
C467 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_557_413# -3.67e-20
C468 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# -0.00466f
C469 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# V_LOW -1.39e-35
C470 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 2.71e-19
C471 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 0.00106f
C472 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 7.96e-20
C473 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.5e-20
C474 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 0.07f
C475 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 0.03f
C476 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_557_413# -0.0012f
C477 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# -0.00641f
C478 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.35e-19
C479 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 9.84e-20
C480 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__nor2_1_0/Y 0.00301f
C481 RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_30/HI 1.89e-19
C482 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_24/HI 0.21f
C483 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_23/LO 6.51e-21
C484 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# -0.00385f
C485 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 1.42e-32
C486 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 2.2e-20
C487 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# -0.00491f
C488 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_891_329# -0.00159f
C489 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# V_LOW -0.0229f
C490 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# 3.75e-21
C491 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 2.19e-19
C492 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 2.19e-19
C493 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0307f
C494 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__conb_1_45/HI 0.0309f
C495 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 5.66e-19
C496 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 5.66e-19
C497 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 5.74e-21
C498 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 5.16e-20
C499 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__conb_1_44/HI 2.5e-21
C500 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 5.66e-20
C501 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__conb_1_47/HI 0.00314f
C502 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_11/LO 9.95e-20
C503 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# -6.57e-19
C504 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__conb_1_36/HI 6.78e-19
C505 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.77e-21
C506 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.78e-22
C507 FULL_COUNTER.COUNT_SUB_DFF11.Q V_LOW 1.41f
C508 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__conb_1_22/HI 1.63e-19
C509 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nand3_1_2/B 1.99e-19
C510 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.00191f
C511 sky130_fd_sc_hd__conb_1_42/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0198f
C512 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__inv_1_49/Y 0.0103f
C513 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 6.82e-19
C514 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/Q_N -8.88e-34
C515 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 0.0135f
C516 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 6.31e-21
C517 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 3.23e-21
C518 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# V_LOW -0.00121f
C519 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 3.05e-19
C520 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 7.14e-20
C521 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# V_LOW 1.79e-20
C522 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 1.15e-19
C523 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# V_GND -0.0041f
C524 sky130_fd_sc_hd__dfbbn_1_40/Q_N V_LOW -0.00509f
C525 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_13/LO 1.03e-19
C526 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_5/HI 7.91e-20
C527 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0013f
C528 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# V_LOW -1.39e-35
C529 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# V_GND 0.0136f
C530 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__inv_1_15/Y 0.00152f
C531 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__conb_1_2/LO 7.93e-21
C532 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# 4.17e-19
C533 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# V_GND 0.00549f
C534 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 2.45e-20
C535 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0.00592f
C536 sky130_fd_sc_hd__inv_1_109/Y FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.85e-20
C537 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0.00592f
C538 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 2.45e-20
C539 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 1.91e-19
C540 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 5.95e-19
C541 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_19/LO 1.53e-19
C542 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__inv_1_15/Y 5.4e-19
C543 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 3.28e-20
C544 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 1.4e-21
C545 RISING_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 3.52e-20
C546 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 0.00113f
C547 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_DFF14.Q 3.03f
C548 sky130_fd_sc_hd__conb_1_26/LO RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0382f
C549 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_103/Y 0.0385f
C550 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00147f
C551 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0366f
C552 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# V_GND 0.00244f
C553 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_1_108/Y 4.4e-19
C554 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# -0.00117f
C555 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# -6.22e-19
C556 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# -0.00811f
C557 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# V_LOW 1.38e-19
C558 sky130_fd_sc_hd__inv_1_90/Y V_LOW 0.371f
C559 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1e-20
C560 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# V_GND -3.83e-19
C561 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 3.55e-20
C562 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_61/Y 0.024f
C563 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__conb_1_28/HI 4.26e-20
C564 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_16_2/Y 2.97e-21
C565 sky130_fd_sc_hd__nand2_1_2/A V_LOW 0.0543f
C566 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.13e-20
C567 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 6.1e-19
C568 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 6.47e-22
C569 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00291f
C570 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00238f
C571 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 4.32e-19
C572 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.1e-21
C573 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 2.59e-21
C574 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00382f
C575 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 4.71e-20
C576 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 2.01e-20
C577 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_23/Y 0.0654f
C578 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 7.69e-20
C579 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_43/A 0.00152f
C580 sky130_fd_sc_hd__inv_1_17/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0247f
C581 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# sky130_fd_sc_hd__conb_1_8/HI 6.95e-21
C582 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__conb_1_5/HI 0.00267f
C583 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.81e-19
C584 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__conb_1_34/HI 7.78e-19
C585 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# V_GND 0.00104f
C586 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# sky130_fd_sc_hd__conb_1_51/HI 3.52e-19
C587 sky130_fd_sc_hd__dfbbn_1_4/Q_N V_LOW -0.00958f
C588 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_32/HI 4.56e-21
C589 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00186f
C590 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 1.71e-20
C591 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 2.97e-19
C592 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 1.99e-20
C593 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 2.27e-19
C594 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 8.79e-21
C595 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 4.81e-21
C596 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 6.25e-19
C597 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.00449f
C598 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_16/HI 3.78e-19
C599 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# V_LOW 1.38e-19
C600 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 2.98e-20
C601 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# 1.81e-20
C602 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__inv_1_12/Y 0.00291f
C603 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.32e-20
C604 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__conb_1_33/LO 2.41e-20
C605 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_19/Y 4.43e-21
C606 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 2.09e-21
C607 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# 7.58e-19
C608 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_23/HI 0.00566f
C609 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.583f
C610 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00497f
C611 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 4.32e-21
C612 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 3.22e-20
C613 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00244f
C614 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 1.38e-20
C615 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# -3.46e-20
C616 sky130_fd_sc_hd__conb_1_3/HI CLOCK_GEN.SR_Op.Q 0.00285f
C617 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__conb_1_2/HI 0.0351f
C618 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# V_LOW -6.55e-19
C619 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# -4.66e-20
C620 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_381_47# -3.79e-20
C621 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 7.8e-21
C622 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_103/Y 0.0366f
C623 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00485f
C624 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__conb_1_47/HI 0.0338f
C625 sky130_fd_sc_hd__dfbbn_1_43/a_557_413# V_LOW 3.56e-20
C626 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# sky130_fd_sc_hd__inv_1_13/Y 3.81e-20
C627 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# sky130_fd_sc_hd__inv_1_8/Y 7.05e-19
C628 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# V_LOW 4.8e-20
C629 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# sky130_fd_sc_hd__conb_1_22/HI 1.99e-21
C630 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# V_GND 9.11e-19
C631 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.87e-20
C632 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_581_47# 1.96e-19
C633 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_193_47# 0.0398f
C634 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__conb_1_3/HI 2.89e-20
C635 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 2.78e-20
C636 sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# V_GND -0.00159f
C637 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 7.98e-19
C638 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 0.00104f
C639 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 1.94e-19
C640 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 3.46e-19
C641 sky130_fd_sc_hd__conb_1_49/LO V_LOW -0.00433f
C642 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0012f
C643 sky130_fd_sc_hd__dfbbn_1_7/Q_N V_LOW -0.00229f
C644 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.0199f
C645 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# V_GND 1.59e-19
C646 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# -0.00155f
C647 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# -0.0152f
C648 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.68e-20
C649 Reset sky130_fd_sc_hd__inv_16_2/Y 0.0705f
C650 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# 2.01e-20
C651 sky130_fd_sc_hd__dfbbn_1_3/a_581_47# V_GND 4.71e-19
C652 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_27_47# 0.0014f
C653 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 2.89e-19
C654 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_791_47# 4e-19
C655 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 4e-19
C656 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 2.89e-19
C657 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__inv_1_15/Y 5.37e-21
C658 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.98e-20
C659 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.112f
C660 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/Q_N -7.69e-20
C661 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 0.0107f
C662 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__inv_1_16/Y 1.31e-20
C663 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__inv_1_108/Y 0.00222f
C664 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# V_GND 0.0404f
C665 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# 8.93e-20
C666 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -6.22e-19
C667 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# -0.00242f
C668 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# -0.00827f
C669 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_40/a_27_47# 0.183f
C670 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_94/A 8.37e-19
C671 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__inv_1_47/Y 3.56e-19
C672 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0.0111f
C673 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF3.Q 3.05e-20
C674 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.03e-20
C675 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.6e-19
C676 sky130_fd_sc_hd__nand2_8_0/a_27_47# V_GND 0.056f
C677 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_1_100/Y 0.0573f
C678 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_41/HI 0.274f
C679 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_16_2/Y 3.83e-19
C680 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 1.29e-20
C681 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00153f
C682 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00155f
C683 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.63e-21
C684 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__conb_1_48/LO 2.72e-20
C685 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.98e-21
C686 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 8.45e-19
C687 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0365f
C688 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.17e-20
C689 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00156f
C690 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__conb_1_5/HI 6.51e-21
C691 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0211f
C692 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00145f
C693 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.11e-19
C694 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 2.81e-20
C695 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 8.08e-21
C696 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 3.16e-19
C697 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 2.69e-19
C698 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 7.55e-19
C699 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00184f
C700 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_21/HI 5.54e-21
C701 sky130_fd_sc_hd__nand2_8_7/a_27_47# V_LOW -0.00286f
C702 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 2.96e-19
C703 FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.18e-20
C704 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 2.38e-20
C705 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.53e-19
C706 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/Q_N 3.21e-19
C707 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__conb_1_33/HI 0.017f
C708 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00285f
C709 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# -0.00344f
C710 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# -6.43e-20
C711 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 1.07e-19
C712 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 3.02e-21
C713 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 8.05e-20
C714 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__conb_1_35/LO 4.55e-20
C715 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 1.75e-20
C716 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_6/HI 9.8e-21
C717 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__inv_1_15/Y 4.06e-19
C718 sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__inv_16_1/Y 1.33e-20
C719 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nand3_1_2/B 1.87e-20
C720 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0368f
C721 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00439f
C722 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_791_47# 0.0037f
C723 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00103f
C724 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# 6.75e-20
C725 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.00112f
C726 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 0.00177f
C727 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_16_2/Y 0.322f
C728 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# V_LOW 0.013f
C729 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# V_LOW 0.00298f
C730 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 0.00154f
C731 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00534f
C732 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# V_LOW 3.56e-20
C733 sky130_fd_sc_hd__inv_1_2/Y V_SENSE 0.0619f
C734 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# V_LOW 0.0161f
C735 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# -1.24e-20
C736 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# 5.22e-19
C737 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 4.93e-20
C738 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.105f
C739 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_19/Y 4.5e-20
C740 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.207f
C741 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# V_LOW -0.0267f
C742 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 1.07e-20
C743 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 0.0093f
C744 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.19e-19
C745 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 9.79e-19
C746 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 3.85e-19
C747 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__inv_16_0/Y 2.27e-21
C748 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# V_LOW 0.0155f
C749 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_50/Y 2.17e-19
C750 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# V_GND -0.00526f
C751 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# V_GND -0.00802f
C752 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# V_LOW 0.0186f
C753 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_22/HI 2.97e-19
C754 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__conb_1_28/LO 4.13e-19
C755 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.0764f
C756 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# -5.77e-20
C757 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# -2.52e-19
C758 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# V_GND 1.69e-19
C759 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0262f
C760 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# V_GND 0.0018f
C761 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/Q_N 9.8e-20
C762 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 0.0074f
C763 sky130_fd_sc_hd__dfbbn_1_49/a_581_47# sky130_fd_sc_hd__inv_1_47/Y 5.8e-19
C764 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# V_GND 0.00133f
C765 sky130_fd_sc_hd__inv_1_50/A V_LOW 0.418f
C766 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# -0.233f
C767 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__conb_1_45/HI 4.36e-19
C768 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.00121f
C769 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_193_47# -0.233f
C770 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 2.85e-21
C771 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 0.00259f
C772 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.06e-21
C773 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__conb_1_49/HI 0.0923f
C774 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# V_GND 0.00179f
C775 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_1_15/Y 6.84e-19
C776 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_1_59/Y 0.0234f
C777 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0117f
C778 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0197f
C779 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# V_GND -0.0348f
C780 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 2.76e-19
C781 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0011f
C782 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0835f
C783 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.25e-20
C784 sky130_fd_sc_hd__nand2_1_1/a_113_47# V_GND 2.83e-20
C785 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 0.00374f
C786 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0206f
C787 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_1_112/Y 4.37e-21
C788 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_4/HI 1.79e-19
C789 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.27e-20
C790 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# V_LOW -0.103f
C791 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# V_GND 0.0405f
C792 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 0.00154f
C793 sky130_fd_sc_hd__conb_1_16/HI sky130_fd_sc_hd__conb_1_17/HI 8.89e-21
C794 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 2.07e-19
C795 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__nand2_8_6/a_27_47# 0.00656f
C796 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.62e-20
C797 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 8.88e-20
C798 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.56e-20
C799 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/Q_N -2.84e-32
C800 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.27e-19
C801 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# -0.00407f
C802 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 9.03e-19
C803 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0524f
C804 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.97e-20
C805 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00171f
C806 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__inv_1_20/Y 7.05e-19
C807 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 8.5e-22
C808 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 1.55e-20
C809 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 1.11e-19
C810 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__inv_1_62/Y 7.02e-19
C811 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# -0.00138f
C812 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# V_GND -0.00522f
C813 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__conb_1_31/HI 3.62e-20
C814 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__inv_1_11/Y 7.25e-19
C815 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 5.15e-20
C816 sky130_fd_sc_hd__inv_1_45/Y V_GND 0.0877f
C817 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.8e-20
C818 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0045f
C819 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_1_99/Y 0.00193f
C820 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00162f
C821 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00737f
C822 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__conb_1_24/HI 1.7e-19
C823 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__conb_1_45/HI 2.43e-19
C824 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# V_LOW 1.79e-20
C825 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__inv_16_2/Y 0.109f
C826 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 2.75e-20
C827 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_1_17/Y 0.0114f
C828 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 2.62e-19
C829 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 7.26e-20
C830 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 4.3e-20
C831 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__conb_1_38/LO 6.57e-20
C832 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_95/A 8.06e-19
C833 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_581_47# -2.6e-20
C834 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 4.39e-19
C835 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00783f
C836 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_9/Y 3.84e-19
C837 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 0.00295f
C838 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# V_LOW 1.79e-20
C839 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 1.6e-19
C840 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__conb_1_0/HI 1.36e-20
C841 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# V_LOW 0.00185f
C842 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00431f
C843 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__inv_16_1/Y 8.37e-19
C844 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# 4.84e-20
C845 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_108/Y 2.73e-19
C846 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_1_58/Y 0.00258f
C847 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.2e-19
C848 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 8.58e-20
C849 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.284f
C850 sky130_fd_sc_hd__conb_1_33/LO V_LOW 0.0408f
C851 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 0.00144f
C852 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 3.76e-20
C853 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 3.76e-20
C854 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 0.00144f
C855 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# V_LOW 1.79e-20
C856 sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF11.Q 3.11e-20
C857 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_1_17/Y 9.84e-20
C858 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# V_GND -3.53e-19
C859 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__inv_1_50/Y 1.64e-21
C860 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# V_GND 0.00277f
C861 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__inv_16_2/Y 0.0557f
C862 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_105/Y 0.00316f
C863 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.207f
C864 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# 0.0351f
C865 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# -1.76e-19
C866 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.335f
C867 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.00475f
C868 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# V_GND -0.00167f
C869 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/Q_N -9.56e-20
C870 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00109f
C871 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_11/HI 0.0455f
C872 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 2.77e-20
C873 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_39/HI 1.68e-19
C874 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# V_GND 1.48e-19
C875 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# V_LOW 3.56e-20
C876 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__inv_1_61/Y 0.00344f
C877 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# CLOCK_GEN.SR_Op.Q 1.75e-19
C878 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 0.00171f
C879 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# V_GND 0.00122f
C880 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.117f
C881 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.00519f
C882 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__conb_1_46/HI 0.00121f
C883 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 1.62e-19
C884 sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00751f
C885 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0239f
C886 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 6.8e-19
C887 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__conb_1_6/HI 0.00239f
C888 sky130_fd_sc_hd__inv_1_55/Y V_GND 0.0144f
C889 FULL_COUNTER.COUNT_SUB_DFF0.Q CLOCK_GEN.SR_Op.Q 6.33e-19
C890 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# sky130_fd_sc_hd__conb_1_49/HI 0.00216f
C891 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand2_8_3/A 0.0607f
C892 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 5.73e-21
C893 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# V_GND -3.53e-19
C894 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__inv_1_15/Y 0.00138f
C895 sky130_fd_sc_hd__dfbbn_1_42/a_581_47# sky130_fd_sc_hd__inv_1_59/Y 6.07e-19
C896 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0352f
C897 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# V_GND 2.94e-19
C898 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 4.85e-19
C899 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00562f
C900 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0195f
C901 sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0021f
C902 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_381_47# 0.00186f
C903 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 0.0275f
C904 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# 5.15e-19
C905 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.167f
C906 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -2.18e-19
C907 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -0.00226f
C908 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 2.13e-32
C909 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# V_GND 1.68e-19
C910 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# V_LOW -9.94e-19
C911 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# -6.29e-19
C912 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_557_413# -3.67e-20
C913 sky130_fd_sc_hd__fill_4_56/VPB V_GND 0.441f
C914 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_5/HI 1.24e-19
C915 sky130_fd_sc_hd__inv_1_100/Y V_GND 0.121f
C916 sky130_fd_sc_hd__conb_1_21/HI sky130_fd_sc_hd__conb_1_17/HI 2.75e-20
C917 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.85e-21
C918 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.94e-19
C919 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 6.62e-20
C920 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -0.0528f
C921 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_581_47# -2.6e-20
C922 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_97/A 4.71e-20
C923 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0648f
C924 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_1_99/Y 1.21e-19
C925 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 0.0242f
C926 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_1_63/Y 1.39e-19
C927 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# -3.86e-20
C928 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# -1.03e-19
C929 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# -9.32e-20
C930 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.3e-19
C931 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# V_GND 1.46e-19
C932 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# sky130_fd_sc_hd__inv_1_11/Y 2.57e-19
C933 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# -0.00263f
C934 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# -0.00226f
C935 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -2.18e-19
C936 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.9e-19
C937 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.013f
C938 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__inv_1_99/Y 0.00599f
C939 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 3.5e-19
C940 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00532f
C941 sky130_fd_sc_hd__inv_1_102/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.138f
C942 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.8e-20
C943 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0244f
C944 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.46e-20
C945 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00396f
C946 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# V_LOW 0.00243f
C947 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 1.8e-21
C948 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# -5.54e-21
C949 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# -1.6e-19
C950 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# -2.6e-19
C951 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.7e-19
C952 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.66e-19
C953 sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__inv_16_1/Y 0.411f
C954 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 1.59e-19
C955 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__conb_1_34/LO 0.0011f
C956 sky130_fd_sc_hd__inv_1_49/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.126f
C957 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_1/LO 0.00375f
C958 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_51/A 0.0494f
C959 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 6.41e-19
C960 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__inv_1_5/Y 1.25e-19
C961 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 5.43e-37
C962 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00873f
C963 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.46e-19
C964 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__inv_1_90/Y 0.00707f
C965 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00237f
C966 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_9/Y 0.0941f
C967 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.47e-21
C968 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# sky130_fd_sc_hd__inv_1_105/Y 9.3e-22
C969 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# V_GND 3.73e-19
C970 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_1_22/Y 0.0747f
C971 sky130_fd_sc_hd__conb_1_42/HI FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0229f
C972 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0727f
C973 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# V_LOW 0.00466f
C974 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_557_413# -3.67e-20
C975 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# -0.00793f
C976 FULL_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 1.28e-20
C977 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 1.06e-19
C978 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_71/A 0.0364f
C979 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.03e-19
C980 sky130_fd_sc_hd__inv_2_0/Y V_SENSE 1.08f
C981 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_37/HI -0.00109f
C982 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# 3.92e-21
C983 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# V_GND -0.00141f
C984 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 2.15e-19
C985 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 6.95e-20
C986 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0.0346f
C987 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0109f
C988 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 5.51e-21
C989 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 1.25e-19
C990 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00292f
C991 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 1.71e-20
C992 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 4.39e-21
C993 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_891_329# -0.00159f
C994 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# -0.00524f
C995 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 8.2e-19
C996 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_1_19/Y 2.43e-20
C997 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_68/A 0.00304f
C998 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# 5.52e-20
C999 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__conb_1_6/HI 0.00343f
C1000 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# sky130_fd_sc_hd__conb_1_42/HI 4.16e-20
C1001 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 2.84e-19
C1002 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 9.41e-19
C1003 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0528f
C1004 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 7.04e-20
C1005 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 3.81e-19
C1006 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# V_GND 9.12e-19
C1007 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# 1.12e-19
C1008 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 3.01e-21
C1009 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00251f
C1010 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 8.84e-20
C1011 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# -2.65e-20
C1012 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_12/HI 2.07e-19
C1013 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__conb_1_40/HI 0.00187f
C1014 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 4.57e-21
C1015 sky130_fd_sc_hd__conb_1_24/HI V_LOW 0.0443f
C1016 sky130_fd_sc_hd__inv_1_109/Y FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.303f
C1017 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 1.66e-20
C1018 sky130_fd_sc_hd__inv_1_0/A V_GND 0.0852f
C1019 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 4.22e-21
C1020 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# -4.66e-20
C1021 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_381_47# -3.79e-20
C1022 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0283f
C1023 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# CLOCK_GEN.SR_Op.Q 1.85e-19
C1024 sky130_fd_sc_hd__inv_1_61/Y V_LOW 0.154f
C1025 sky130_fd_sc_hd__conb_1_7/HI V_LOW 0.18f
C1026 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_41/LO 3.78e-19
C1027 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 7.39e-19
C1028 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# 4.54e-19
C1029 sky130_fd_sc_hd__conb_1_44/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0445f
C1030 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# sky130_fd_sc_hd__inv_1_63/Y 2.07e-21
C1031 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 4.11e-21
C1032 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 5.09e-20
C1033 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 3.13e-19
C1034 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.00382f
C1035 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00128f
C1036 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# -2.57e-20
C1037 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_21/HI 0.0726f
C1038 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0355f
C1039 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/Q_N -4.16e-20
C1040 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.24e-20
C1041 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__conb_1_50/LO 0.0116f
C1042 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# -9.32e-20
C1043 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0024f
C1044 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# V_LOW -0.109f
C1045 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 4.26e-20
C1046 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.66e-20
C1047 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_891_329# 2.44e-19
C1048 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# -9.32e-20
C1049 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 5.54e-19
C1050 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# V_LOW -2.78e-35
C1051 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_53/Y 3.13e-20
C1052 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/Q_N 5.44e-20
C1053 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.22e-19
C1054 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 2.47e-19
C1055 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_8/HI 1.04e-19
C1056 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.0016f
C1057 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 0.0016f
C1058 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__conb_1_6/HI 5.93e-19
C1059 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__nand3_1_0/Y 3.33e-19
C1060 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 6.4e-20
C1061 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 1.44e-19
C1062 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 6.4e-19
C1063 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.06e-21
C1064 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.01e-22
C1065 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.00322f
C1066 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.9e-20
C1067 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__conb_1_48/HI 3.32e-19
C1068 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.00178f
C1069 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__inv_1_16/Y 0.00634f
C1070 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# V_GND -0.00489f
C1071 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_93/A 1.44e-20
C1072 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0446f
C1073 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0175f
C1074 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_31/HI 1.51e-19
C1075 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 7.04e-19
C1076 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 0.0115f
C1077 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.17e-19
C1078 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# 6.45e-19
C1079 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.35e-20
C1080 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__conb_1_24/HI 4.06e-20
C1081 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# V_GND 0.00825f
C1082 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 1.73e-20
C1083 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00694f
C1084 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# -0.00385f
C1085 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_97/Y 7.6e-19
C1086 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__inv_1_19/Y 1.33e-21
C1087 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_108/Y 8.99e-21
C1088 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__conb_1_17/HI 8.11e-21
C1089 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__conb_1_42/HI 0.00713f
C1090 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0197f
C1091 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__conb_1_27/HI 1.33e-19
C1092 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/Q_N -4.33e-20
C1093 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.47e-20
C1094 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__conb_1_40/HI 0.00586f
C1095 FALLING_COUNTER.COUNT_SUB_DFF2.Q V_GND 0.586f
C1096 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.54e-20
C1097 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__inv_1_93/A 4.29e-20
C1098 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 3.99e-19
C1099 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_1_8/Y 1.23e-19
C1100 sky130_fd_sc_hd__dfbbn_1_5/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00373f
C1101 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__conb_1_7/LO 4.01e-21
C1102 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__inv_1_56/Y 0.00605f
C1103 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_39/Q_N 1.19e-20
C1104 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_55/Y 5.77e-19
C1105 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__conb_1_34/LO 6.57e-20
C1106 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_32/Y 0.0443f
C1107 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1_1/Y 4.68e-20
C1108 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y 0.14f
C1109 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/A 0.183f
C1110 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 1.72e-19
C1111 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__conb_1_23/HI -0.0541f
C1112 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/Q_N -4.33e-20
C1113 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.0299f
C1114 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 5.67e-21
C1115 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 5.25e-19
C1116 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 6.25e-19
C1117 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# V_LOW -9.94e-19
C1118 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# 5.86e-21
C1119 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_12/HI 7.7e-21
C1120 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0.00811f
C1121 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__conb_1_3/LO 0.0209f
C1122 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.57e-20
C1123 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/Q_N -4.33e-20
C1124 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_25/HI -8.83e-19
C1125 sky130_fd_sc_hd__dfbbn_1_30/Q_N V_LOW -9.22e-19
C1126 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00162f
C1127 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.32e-20
C1128 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__conb_1_2/HI 0.00128f
C1129 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 1.03e-19
C1130 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_76/A 0.00113f
C1131 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# 0.00412f
C1132 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.68e-19
C1133 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_101/Y -1.12e-19
C1134 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.03e-19
C1135 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_791_47# 7.41e-19
C1136 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 4.18e-19
C1137 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00133f
C1138 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_21/Y 8.87e-19
C1139 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_38/LO 5.49e-19
C1140 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# V_LOW -0.00266f
C1141 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# CLOCK_GEN.SR_Op.Q 0.0061f
C1142 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_42/Y 0.0183f
C1143 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 1.64e-20
C1144 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__conb_1_12/HI 5.44e-19
C1145 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 7.66e-21
C1146 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF3.Q 5.47e-21
C1147 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# V_GND 1.59e-19
C1148 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__inv_1_54/Y 1.72e-20
C1149 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 2.19e-19
C1150 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_75/A 0.00747f
C1151 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.94e-20
C1152 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 6.4e-19
C1153 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.15e-19
C1154 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00596f
C1155 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 9.49e-19
C1156 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00378f
C1157 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__conb_1_51/HI 6.92e-19
C1158 sky130_fd_sc_hd__dfbbn_1_35/Q_N V_LOW -0.00509f
C1159 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__inv_1_11/Y 2.16e-20
C1160 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__conb_1_39/HI 0.00101f
C1161 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0232f
C1162 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 5.13e-19
C1163 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_40/HI 0.00125f
C1164 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__inv_1_18/Y 2.92e-19
C1165 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.0018f
C1166 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 5.09e-21
C1167 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# sky130_fd_sc_hd__conb_1_24/HI 5.18e-21
C1168 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# V_GND 4.43e-19
C1169 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__conb_1_6/HI 0.00163f
C1170 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/Q_N -6.48e-19
C1171 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_92/Y 0.00424f
C1172 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 1.18e-19
C1173 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 3.87e-19
C1174 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0155f
C1175 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 0.0259f
C1176 sky130_fd_sc_hd__conb_1_18/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 9.35e-20
C1177 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0.00609f
C1178 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# CLOCK_GEN.SR_Op.Q 4.7e-20
C1179 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__conb_1_22/HI 0.00135f
C1180 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00111f
C1181 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_11/HI 2.5e-20
C1182 sky130_fd_sc_hd__conb_1_1/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0143f
C1183 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# V_LOW 0.0688f
C1184 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_49/HI 0.0216f
C1185 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_891_329# 0.00134f
C1186 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# V_GND 0.00443f
C1187 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 1.28e-20
C1188 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.68e-19
C1189 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.89e-19
C1190 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00308f
C1191 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__inv_1_99/Y 8.09e-19
C1192 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 7.98e-20
C1193 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# sky130_fd_sc_hd__conb_1_21/HI 0.00211f
C1194 RISING_COUNTER.COUNT_SUB_DFF0.Q CLOCK_GEN.SR_Op.Q 0.451f
C1195 sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 3.37e-19
C1196 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_43/Y 6.57e-19
C1197 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__inv_1_19/Y 0.00563f
C1198 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.00613f
C1199 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_50/a_473_413# 4.15e-20
C1200 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_381_47# 7.43e-20
C1201 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# -0.00222f
C1202 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# -7.6e-19
C1203 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_30/HI 1.09e-19
C1204 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# -3.48e-20
C1205 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_891_329# -2.2e-20
C1206 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 8.03e-21
C1207 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__inv_1_6/Y 8.46e-19
C1208 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_43/Q_N -2.84e-32
C1209 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 3.72e-19
C1210 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.09e-21
C1211 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0156f
C1212 sky130_fd_sc_hd__inv_1_119/Y V_GND 0.498f
C1213 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# V_GND 0.00834f
C1214 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_18/HI 0.108f
C1215 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# V_GND 0.00729f
C1216 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 4.26e-21
C1217 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# sky130_fd_sc_hd__inv_1_58/Y 1.19e-19
C1218 sky130_fd_sc_hd__conb_1_37/HI V_LOW 0.169f
C1219 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_13/Q_N 1.01e-19
C1220 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 0.00516f
C1221 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# V_GND 0.00929f
C1222 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_791_47# 4.35e-20
C1223 sky130_fd_sc_hd__conb_1_50/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.145f
C1224 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0.00526f
C1225 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 0.019f
C1226 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# sky130_fd_sc_hd__conb_1_12/HI 9.94e-22
C1227 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_28/HI -0.00351f
C1228 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 0.00554f
C1229 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00197f
C1230 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_106/Y 0.0622f
C1231 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/Q_N 0.0248f
C1232 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.86e-20
C1233 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# -0.0147f
C1234 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_647_21# -6.43e-20
C1235 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_6/HI 0.23f
C1236 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 1.27e-19
C1237 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_891_329# 0.00186f
C1238 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_12/HI 0.00854f
C1239 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_24/a_791_47# 5.13e-19
C1240 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.78e-19
C1241 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# -3.79e-20
C1242 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# -4.66e-20
C1243 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__conb_1_37/HI 1.79e-19
C1244 sky130_fd_sc_hd__conb_1_49/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.38e-19
C1245 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 1.83e-20
C1246 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 0.188f
C1247 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 9.97e-19
C1248 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 3.55e-21
C1249 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 2.84e-20
C1250 FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 1.66f
C1251 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__conb_1_22/HI 2.5e-19
C1252 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# -0.00312f
C1253 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# -0.00746f
C1254 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.108f
C1255 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.35e-20
C1256 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_13/Y 0.0913f
C1257 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__inv_1_18/Y 1.02e-19
C1258 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__conb_1_16/HI 0.0015f
C1259 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.72e-21
C1260 sky130_fd_sc_hd__dfbbn_1_28/Q_N RISING_COUNTER.COUNT_SUB_DFF3.Q 1.83e-19
C1261 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 9.94e-20
C1262 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.25e-20
C1263 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# V_LOW 4.8e-20
C1264 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.55e-19
C1265 sky130_fd_sc_hd__inv_1_14/Y V_GND 0.258f
C1266 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# V_LOW 0.014f
C1267 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_941_21# 4.88e-20
C1268 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_5/Y 0.0538f
C1269 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_16_1/Y 0.00178f
C1270 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_75/A 0.124f
C1271 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__conb_1_12/HI -5.67e-19
C1272 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 2.44e-20
C1273 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 2.94e-19
C1274 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 1.5e-20
C1275 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__inv_1_102/Y 2.39e-19
C1276 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# V_LOW -0.00477f
C1277 sky130_fd_sc_hd__inv_1_93/A V_LOW 0.26f
C1278 sky130_fd_sc_hd__dfbbn_1_7/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00163f
C1279 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# -4.1e-19
C1280 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_891_329# -2.2e-20
C1281 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_1_15/Y 0.0137f
C1282 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.41e-19
C1283 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 5.49e-20
C1284 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 8.86e-22
C1285 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 9.16e-20
C1286 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__conb_1_6/HI -2.07e-19
C1287 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# V_GND -0.174f
C1288 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.53e-20
C1289 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.36e-19
C1290 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 2.2e-20
C1291 FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_107/Y 0.329f
C1292 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_791_47# 5.14e-19
C1293 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 7.89e-20
C1294 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_18/Y 0.0969f
C1295 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 1.31e-20
C1296 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# -0.00591f
C1297 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# -6.43e-20
C1298 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 8.5e-21
C1299 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# V_LOW 2.94e-20
C1300 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_1_57/Y 4.19e-19
C1301 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# V_GND 1.47e-19
C1302 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_65/Y 2.16e-21
C1303 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand2_8_9/Y 0.00624f
C1304 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 0.02f
C1305 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# V_GND 0.00324f
C1306 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00265f
C1307 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.91e-20
C1308 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__inv_1_99/Y -2.87e-20
C1309 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.109f
C1310 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# V_LOW 2.26e-20
C1311 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 8.78e-21
C1312 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0338f
C1313 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00422f
C1314 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 2.76e-21
C1315 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# V_LOW 2.26e-20
C1316 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__conb_1_35/HI 0.0399f
C1317 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# V_GND 2.27e-19
C1318 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.62e-21
C1319 sky130_fd_sc_hd__conb_1_22/LO V_GND -0.00146f
C1320 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 3.21e-20
C1321 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 3.1e-20
C1322 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__inv_16_2/Y 0.909f
C1323 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 2.7e-20
C1324 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 9.06e-19
C1325 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__conb_1_40/HI 0.00633f
C1326 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 5.62e-19
C1327 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 4.08e-19
C1328 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 2.64e-19
C1329 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 7e-19
C1330 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 9.33e-19
C1331 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00391f
C1332 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0139f
C1333 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__conb_1_9/HI 3.5e-22
C1334 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# -9.32e-20
C1335 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# -0.00142f
C1336 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__conb_1_42/HI 1.36e-19
C1337 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 1.04e-19
C1338 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_1_103/Y 0.00105f
C1339 sky130_fd_sc_hd__inv_1_46/Y V_LOW 0.163f
C1340 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00415f
C1341 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.05f
C1342 sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# V_GND 0.00144f
C1343 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_63/Y 3.43e-19
C1344 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__nand3_1_0/Y 0.00209f
C1345 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# V_GND 0.00172f
C1346 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__conb_1_38/HI 0.0191f
C1347 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# V_LOW 0.00576f
C1348 sky130_fd_sc_hd__inv_1_111/Y RISING_COUNTER.COUNT_SUB_DFF1.Q 9.78e-20
C1349 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# V_GND 0.00306f
C1350 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00278f
C1351 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# V_LOW -0.00118f
C1352 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 9.71e-19
C1353 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 3.15e-19
C1354 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 0.00342f
C1355 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 7.08e-20
C1356 sky130_fd_sc_hd__inv_1_71/A CLOCK_GEN.SR_Op.Q 6.97e-19
C1357 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 1.11e-20
C1358 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 1.1e-19
C1359 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_76/A 0.00101f
C1360 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_9/LO 0.00125f
C1361 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__conb_1_33/HI 0.00126f
C1362 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.523f
C1363 sky130_fd_sc_hd__inv_1_10/Y V_LOW 0.424f
C1364 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# -0.0144f
C1365 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_891_329# -0.00159f
C1366 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__inv_16_1/Y 2.81e-20
C1367 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_21/HI 1.18e-20
C1368 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 6.26e-20
C1369 sky130_fd_sc_hd__dfbbn_1_28/Q_N RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00671f
C1370 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__conb_1_12/HI 0.0239f
C1371 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 9.39e-22
C1372 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_83/Y 0.1f
C1373 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__conb_1_26/HI 4.95e-19
C1374 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# -3.48e-20
C1375 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_891_329# -2.2e-20
C1376 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# V_LOW -9.15e-19
C1377 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# 0.00211f
C1378 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# V_GND 4.23e-19
C1379 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_75/A 0.99f
C1380 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__conb_1_22/HI 4.32e-20
C1381 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# V_GND 3.26e-19
C1382 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__conb_1_16/HI 0.00126f
C1383 sky130_fd_sc_hd__nand3_1_1/a_193_47# V_LOW -4.69e-19
C1384 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.78e-19
C1385 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_85/A 1.02e-19
C1386 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# V_LOW 1.79e-20
C1387 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# sky130_fd_sc_hd__conb_1_12/HI -0.00127f
C1388 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# -0.0109f
C1389 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# -6.43e-20
C1390 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_17/HI 1.27e-19
C1391 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.0247f
C1392 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_40/HI 0.00621f
C1393 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 9.83e-21
C1394 sky130_fd_sc_hd__nand3_1_0/Y Reset 0.116f
C1395 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# V_LOW 2.04e-19
C1396 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 1.42e-32
C1397 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# -0.00385f
C1398 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 8.74e-21
C1399 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0075f
C1400 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.71e-19
C1401 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0321f
C1402 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# V_GND 1.2e-19
C1403 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.01e-20
C1404 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0145f
C1405 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.31e-20
C1406 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 1.38e-20
C1407 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 9.03e-20
C1408 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 5.86e-19
C1409 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 0.00327f
C1410 sky130_fd_sc_hd__inv_1_111/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 6.79e-20
C1411 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 5.22e-21
C1412 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0522f
C1413 FULL_COUNTER.COUNT_SUB_DFF15.Q V_LOW 4.5f
C1414 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# sky130_fd_sc_hd__inv_1_18/Y 0.00175f
C1415 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_791_47# 0.00838f
C1416 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00539f
C1417 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__inv_1_57/Y 4.07e-20
C1418 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_13/HI 0.00787f
C1419 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# V_GND 0.0355f
C1420 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# sky130_fd_sc_hd__inv_16_1/Y 0.00113f
C1421 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# V_GND 1.89e-19
C1422 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# -0.00144f
C1423 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0663f
C1424 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0307f
C1425 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.024f
C1426 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_1_99/Y 0.00772f
C1427 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__conb_1_32/HI 0.0288f
C1428 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.121f
C1429 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.46e-20
C1430 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__conb_1_35/HI 9.26e-20
C1431 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_12/LO 0.00869f
C1432 sky130_fd_sc_hd__inv_1_98/Y V_GND 0.103f
C1433 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# -2.01e-20
C1434 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# -0.00263f
C1435 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# Reset 1.17e-19
C1436 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 5.36e-20
C1437 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 1.19e-19
C1438 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_3/LO 0.0652f
C1439 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__conb_1_40/HI 8.88e-20
C1440 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.49e-21
C1441 sky130_fd_sc_hd__dfbbn_1_26/a_581_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00184f
C1442 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__conb_1_27/LO 1.71e-19
C1443 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/Q_N -4.24e-20
C1444 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/Q_N -6.48e-19
C1445 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.35e-19
C1446 sky130_fd_sc_hd__dfbbn_1_22/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00857f
C1447 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_58/Y 0.0288f
C1448 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00773f
C1449 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 4.44e-20
C1450 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__conb_1_35/HI 5.8e-21
C1451 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 1.18e-20
C1452 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_23/Y 1.68e-19
C1453 FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0831f
C1454 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__conb_1_40/HI 0.00333f
C1455 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# sky130_fd_sc_hd__conb_1_38/HI 3.98e-19
C1456 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# V_LOW 1.26e-20
C1457 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# V_GND 0.0276f
C1458 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00213f
C1459 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# V_GND -3.52e-19
C1460 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 8.54e-19
C1461 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 8.24e-19
C1462 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__inv_1_7/Y 1.72e-19
C1463 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_94/Y 0.00235f
C1464 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.77e-20
C1465 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_43/A 4.48e-20
C1466 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_22/a_647_21# 2.07e-21
C1467 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# -0.00592f
C1468 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 5.15e-21
C1469 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 8.13e-20
C1470 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__conb_1_21/HI 1.5e-20
C1471 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# -0.00497f
C1472 sky130_fd_sc_hd__inv_1_3/A V_SENSE 0.157f
C1473 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# -3.46e-20
C1474 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00101f
C1475 sky130_fd_sc_hd__inv_1_94/A V_LOW 0.992f
C1476 sky130_fd_sc_hd__conb_1_44/LO FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00105f
C1477 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0.0724f
C1478 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_48/HI -0.00183f
C1479 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_55/Y 3.55e-19
C1480 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_58/Y 0.0712f
C1481 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__conb_1_26/HI 3.9e-19
C1482 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__conb_1_46/LO 0.00206f
C1483 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__conb_1_12/HI 0.0129f
C1484 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# V_LOW -7.04e-19
C1485 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# V_LOW 3.56e-20
C1486 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0.00127f
C1487 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 8.32e-19
C1488 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 2.53e-19
C1489 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 0.0149f
C1490 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_1_57/Y 0.0352f
C1491 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# sky130_fd_sc_hd__conb_1_40/HI 1.01e-19
C1492 sky130_fd_sc_hd__dfbbn_1_23/Q_N V_LOW -0.00949f
C1493 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 0.0398f
C1494 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 3.59e-20
C1495 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 3.59e-20
C1496 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 3.17e-19
C1497 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 3.17e-19
C1498 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 9.25e-19
C1499 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_381_47# 0.0165f
C1500 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__inv_1_76/A 1.53e-21
C1501 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0035f
C1502 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00229f
C1503 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0144f
C1504 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 1.42e-19
C1505 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 0.00106f
C1506 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.273f
C1507 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 6.06e-19
C1508 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00286f
C1509 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 0.0826f
C1510 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 9.04e-20
C1511 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# V_GND 3.73e-19
C1512 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# V_GND 1.82e-19
C1513 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# -1.44e-20
C1514 sky130_fd_sc_hd__dfbbn_1_0/Q_N FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00313f
C1515 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# V_LOW 3.56e-20
C1516 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# sky130_fd_sc_hd__conb_1_32/HI 4.8e-19
C1517 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_193_47# 0.0316f
C1518 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__inv_1_112/Y 0.0112f
C1519 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__conb_1_12/LO 0.00169f
C1520 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0354f
C1521 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# -9.32e-20
C1522 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__nand3_1_2/Y 0.0407f
C1523 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__conb_1_40/HI 7.43e-21
C1524 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__nand3_1_0/Y 3.26e-20
C1525 sky130_fd_sc_hd__inv_1_23/Y sky130_fd_sc_hd__conb_1_16/HI 0.0221f
C1526 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF9.Q 0.394f
C1527 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__inv_1_58/Y 0.00222f
C1528 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# -3.79e-20
C1529 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# -4.66e-20
C1530 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0122f
C1531 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# Reset 4.55e-21
C1532 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# Reset 2.14e-19
C1533 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nand2_8_1/a_27_47# 0.0361f
C1534 sky130_fd_sc_hd__dfbbn_1_27/Q_N V_LOW -0.00461f
C1535 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# CLOCK_GEN.SR_Op.Q 8.11e-21
C1536 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_95/A 0.00855f
C1537 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# V_GND 1.42e-19
C1538 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 1.23e-19
C1539 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__conb_1_34/HI 0.0303f
C1540 sky130_fd_sc_hd__dfbbn_1_45/Q_N FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0121f
C1541 sky130_fd_sc_hd__dfbbn_1_47/Q_N V_LOW -0.0101f
C1542 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0259f
C1543 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# -1.66e-19
C1544 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__inv_1_62/Y 1.42e-20
C1545 sky130_fd_sc_hd__inv_1_104/Y V_GND 0.133f
C1546 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__conb_1_11/HI 7.47e-19
C1547 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 2.76e-19
C1548 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_97/A 1.1e-19
C1549 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 5.85e-20
C1550 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_381_47# -0.00367f
C1551 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -6.22e-19
C1552 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -0.00242f
C1553 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 8.84e-21
C1554 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_22/LO 0.00534f
C1555 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.41e-19
C1556 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# -0.00141f
C1557 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_9/HI 3.47e-19
C1558 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 8.1e-19
C1559 sky130_fd_sc_hd__conb_1_1/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00761f
C1560 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__inv_1_112/Y 1.06e-19
C1561 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_791_47# 0.00173f
C1562 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 0.00155f
C1563 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__conb_1_48/HI 2.37e-19
C1564 sky130_fd_sc_hd__inv_1_92/Y V_LOW 0.0927f
C1565 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0.00223f
C1566 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_15/HI 0.0492f
C1567 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# -9.13e-21
C1568 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_891_329# -0.00159f
C1569 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_1_108/Y 3.43e-20
C1570 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# V_LOW 7.13e-20
C1571 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0491f
C1572 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_68/A 0.00539f
C1573 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_70/A 0.00134f
C1574 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_2_0/Y 0.0191f
C1575 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# V_LOW -1.39e-35
C1576 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# 4.85e-20
C1577 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 1.8e-20
C1578 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# sky130_fd_sc_hd__inv_16_1/Y 0.00471f
C1579 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 2.31e-21
C1580 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 2.31e-21
C1581 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__conb_1_5/HI 0.0127f
C1582 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 7.32e-20
C1583 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_16_0/Y 0.293f
C1584 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0223f
C1585 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 0.014f
C1586 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.006f
C1587 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.0108f
C1588 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 8.69e-19
C1589 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__conb_1_26/HI 1.23e-20
C1590 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# V_LOW -0.313f
C1591 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_71/A 2.6e-20
C1592 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__inv_1_71/Y 0.00146f
C1593 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# V_LOW 1.45e-19
C1594 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00202f
C1595 sky130_fd_sc_hd__conb_1_10/LO V_GND -0.0043f
C1596 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_4/HI 0.00434f
C1597 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_70/A 1.47e-19
C1598 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_6/HI 9.71e-21
C1599 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 3.54e-21
C1600 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 6.24e-19
C1601 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# V_GND 3.53e-19
C1602 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 0.0113f
C1603 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 8.77e-20
C1604 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 5.27e-20
C1605 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 0.00174f
C1606 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 0.0291f
C1607 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_61/Y 0.00503f
C1608 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_8_3/A 1.08e-19
C1609 sky130_fd_sc_hd__conb_1_48/LO FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00967f
C1610 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_791_47# 0.00264f
C1611 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0398f
C1612 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_105/Y 3.61e-21
C1613 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/Q_N -4.33e-20
C1614 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.73e-20
C1615 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_71/Y 8.67e-19
C1616 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 6.93e-19
C1617 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 0.171f
C1618 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__conb_1_31/HI 0.0421f
C1619 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# V_GND -0.0457f
C1620 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_69/Y 0.0709f
C1621 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__conb_1_0/HI 0.00286f
C1622 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__conb_1_1/HI -4.53e-19
C1623 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# V_GND 9.17e-19
C1624 sky130_fd_sc_hd__inv_1_48/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0399f
C1625 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# sky130_fd_sc_hd__inv_1_103/Y 3.88e-19
C1626 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__conb_1_36/HI 0.0206f
C1627 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF11.Q 3.97e-19
C1628 sky130_fd_sc_hd__conb_1_2/HI sky130_fd_sc_hd__inv_1_5/Y 0.00221f
C1629 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.77e-19
C1630 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__conb_1_12/LO 1.2e-19
C1631 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_17/LO 4.91e-19
C1632 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__inv_1_61/Y 3.75e-21
C1633 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_16_2/Y 0.138f
C1634 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_78/A 2.24e-19
C1635 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__conb_1_11/HI 0.0113f
C1636 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# sky130_fd_sc_hd__conb_1_34/HI 5.96e-19
C1637 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00155f
C1638 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0061f
C1639 sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__inv_1_101/Y 0.00628f
C1640 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__conb_1_42/HI 0.0124f
C1641 sky130_fd_sc_hd__conb_1_47/HI V_GND 0.294f
C1642 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__conb_1_45/HI 0.00212f
C1643 sky130_fd_sc_hd__inv_1_48/Y V_LOW 0.222f
C1644 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_26/Q_N 8.28e-19
C1645 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0876f
C1646 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI 6.89e-20
C1647 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_19/Y 0.0148f
C1648 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# CLOCK_GEN.SR_Op.Q 1.17e-19
C1649 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__conb_1_11/HI 9.48e-21
C1650 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__conb_1_24/HI 1.57e-20
C1651 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 0.0209f
C1652 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 5.91e-19
C1653 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.38e-19
C1654 sky130_fd_sc_hd__inv_1_22/Y V_GND 0.0255f
C1655 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0261f
C1656 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.85e-21
C1657 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# -1.42e-32
C1658 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# -0.00393f
C1659 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# -0.00216f
C1660 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_1_102/Y 1.31e-19
C1661 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# sky130_fd_sc_hd__conb_1_9/HI 4.95e-19
C1662 sky130_fd_sc_hd__dfbbn_1_19/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.95e-19
C1663 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 1.33e-19
C1664 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_1_56/Y 6.69e-20
C1665 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 4.95e-19
C1666 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 8.12e-22
C1667 sky130_fd_sc_hd__conb_1_0/LO V_GND -0.00255f
C1668 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__inv_1_108/Y 3.37e-19
C1669 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 3.14e-19
C1670 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__conb_1_35/LO 0.0712f
C1671 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_105/Y 5.08e-21
C1672 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 3.14e-20
C1673 sky130_fd_sc_hd__dfbbn_1_17/a_557_413# sky130_fd_sc_hd__inv_1_4/Y 8.17e-19
C1674 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__conb_1_5/LO 1.61e-20
C1675 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 5.22e-19
C1676 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 1.71e-19
C1677 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 1.01e-19
C1678 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 3.72e-21
C1679 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# V_LOW -1.39e-35
C1680 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# -3.46e-20
C1681 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 1.42e-32
C1682 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 2.47e-21
C1683 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 5.13e-21
C1684 sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.59e-19
C1685 sky130_fd_sc_hd__dfbbn_1_33/Q_N V_LOW -0.00141f
C1686 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.05e-20
C1687 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.325f
C1688 sky130_fd_sc_hd__inv_1_6/Y V_GND 0.035f
C1689 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_57/Y 0.173f
C1690 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_75/A 1.97e-19
C1691 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_35/HI 0.262f
C1692 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_94/Y 2.62e-19
C1693 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 0.283f
C1694 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.35e-20
C1695 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.5e-19
C1696 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 3.12e-19
C1697 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__conb_1_29/LO 0.0377f
C1698 sky130_fd_sc_hd__nand2_1_0/Y V_GND 0.17f
C1699 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# 4.98e-19
C1700 sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__conb_1_32/HI 0.0074f
C1701 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 1.69e-19
C1702 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 7.23e-20
C1703 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 4.51e-21
C1704 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 9.57e-19
C1705 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 5.19e-20
C1706 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 1.99e-19
C1707 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 9.03e-21
C1708 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__conb_1_42/HI 0.0207f
C1709 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__conb_1_4/HI 9.37e-21
C1710 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0303f
C1711 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_22/a_941_21# 1.34e-20
C1712 sky130_fd_sc_hd__inv_1_43/Y V_GND 0.076f
C1713 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__conb_1_38/HI 8.19e-21
C1714 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# V_LOW 0.00926f
C1715 sky130_fd_sc_hd__dfbbn_1_9/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0193f
C1716 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.68e-19
C1717 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# 0.0223f
C1718 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 9.02e-19
C1719 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0666f
C1720 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__conb_1_10/HI -0.00581f
C1721 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_791_47# 0.0049f
C1722 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# V_LOW -0.00372f
C1723 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.45e-19
C1724 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# sky130_fd_sc_hd__conb_1_31/HI 4.88e-19
C1725 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# V_GND 1.95e-19
C1726 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__conb_1_9/HI 6.14e-19
C1727 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# -0.00125f
C1728 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# -0.00139f
C1729 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__conb_1_36/HI 0.00217f
C1730 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# sky130_fd_sc_hd__conb_1_1/HI -9.78e-19
C1731 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.97e-20
C1732 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__conb_1_36/HI 0.00631f
C1733 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__conb_1_49/LO 4.61e-19
C1734 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__inv_1_22/Y 2.33e-21
C1735 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 3.08e-19
C1736 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.33e-19
C1737 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_941_21# 2.55e-19
C1738 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 1.92e-20
C1739 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__conb_1_21/HI 2.19e-20
C1740 sky130_fd_sc_hd__inv_1_63/Y sky130_fd_sc_hd__inv_16_2/Y 2.07e-19
C1741 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 0.0142f
C1742 FULL_COUNTER.COUNT_SUB_DFF3.Q Reset 3.1e-19
C1743 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# V_LOW 0.00598f
C1744 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_42/Y 5.04e-20
C1745 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# V_GND 0.0124f
C1746 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# V_LOW 0.0243f
C1747 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# V_LOW 0.0148f
C1748 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0408f
C1749 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# V_GND -0.152f
C1750 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 4.03e-21
C1751 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__conb_1_5/LO 6.28e-20
C1752 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.3e-19
C1753 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__conb_1_32/HI 8.24e-20
C1754 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__conb_1_13/HI 0.00645f
C1755 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__inv_1_10/Y 1.72e-20
C1756 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# V_GND -0.00228f
C1757 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# sky130_fd_sc_hd__conb_1_24/HI -2.65e-20
C1758 sky130_fd_sc_hd__dfbbn_1_18/Q_N FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00615f
C1759 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# 0.00111f
C1760 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 4.66e-19
C1761 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_30/HI 3.28e-21
C1762 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 2.29e-19
C1763 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/Q_N -9.56e-20
C1764 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 3.7e-20
C1765 sky130_fd_sc_hd__conb_1_27/LO RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0173f
C1766 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.00305f
C1767 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0371f
C1768 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.89e-19
C1769 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 2.15e-19
C1770 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0.00103f
C1771 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.95e-21
C1772 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00609f
C1773 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 8.58e-19
C1774 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# V_GND 0.0101f
C1775 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.07e-22
C1776 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# V_GND 0.00631f
C1777 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.23e-19
C1778 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# V_GND -0.00661f
C1779 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__inv_1_112/Y 6.94e-20
C1780 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# sky130_fd_sc_hd__inv_1_21/Y 0.00108f
C1781 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.37e-19
C1782 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0416f
C1783 sky130_fd_sc_hd__dfbbn_1_28/Q_N V_LOW -0.00497f
C1784 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# sky130_fd_sc_hd__inv_1_20/Y 8.48e-20
C1785 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 3.72e-19
C1786 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# V_LOW -0.00324f
C1787 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_53/Y 0.00134f
C1788 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 2.2e-20
C1789 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__inv_1_107/Y 4.54e-20
C1790 sky130_fd_sc_hd__inv_1_18/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 0.032f
C1791 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0246f
C1792 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# -4.5e-20
C1793 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -6.23e-21
C1794 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# 0.00253f
C1795 sky130_fd_sc_hd__inv_1_64/A RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00694f
C1796 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.41e-19
C1797 sky130_fd_sc_hd__conb_1_27/HI CLOCK_GEN.SR_Op.Q 1.23e-19
C1798 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0.0113f
C1799 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 2.03e-20
C1800 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_62/Y 1.54e-20
C1801 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 9.14e-19
C1802 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 7.34e-19
C1803 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 1e-19
C1804 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__conb_1_34/HI 1.98e-20
C1805 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 3.16e-21
C1806 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/Q_N 3.16e-21
C1807 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# V_GND 0.0552f
C1808 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0401f
C1809 FULL_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.03f
C1810 sky130_fd_sc_hd__conb_1_11/HI sky130_fd_sc_hd__inv_1_23/Y 6.3e-19
C1811 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# 5.5e-22
C1812 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 1.18e-20
C1813 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 1.96e-19
C1814 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# 5.81e-20
C1815 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 8.7e-21
C1816 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# V_GND 0.0112f
C1817 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# V_GND -0.00456f
C1818 sky130_fd_sc_hd__conb_1_20/LO V_LOW 0.0823f
C1819 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# -0.00336f
C1820 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_45/HI 0.0322f
C1821 sky130_fd_sc_hd__conb_1_44/HI V_GND -0.179f
C1822 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.79e-21
C1823 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_12/HI 1.29e-21
C1824 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# V_LOW 0.00382f
C1825 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# 0.00542f
C1826 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.00812f
C1827 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_1_60/Y 0.0107f
C1828 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00183f
C1829 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# V_LOW -9.15e-19
C1830 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__conb_1_44/LO 1.58e-20
C1831 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_95/Y 0.00232f
C1832 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_65/Y 5.92e-19
C1833 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__conb_1_9/HI -0.00746f
C1834 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__inv_16_2/Y 0.00603f
C1835 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_16_1/Y 0.258f
C1836 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__conb_1_36/HI 7.31e-19
C1837 V_GND RISING_COUNTER.COUNT_SUB_DFF4.Q 1.99f
C1838 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# V_LOW 3.14e-19
C1839 sky130_fd_sc_hd__inv_1_67/Y V_LOW 1.16f
C1840 sky130_fd_sc_hd__conb_1_13/LO V_LOW 0.0885f
C1841 sky130_fd_sc_hd__dfbbn_1_39/Q_N FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.09e-20
C1842 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_70/A 0.101f
C1843 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.15e-19
C1844 sky130_fd_sc_hd__fill_8_819/VPB V_LOW 0.797f
C1845 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_13/HI 0.0013f
C1846 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_1_101/Y 0.0136f
C1847 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_100/Y 0.0067f
C1848 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# V_GND 6.85e-19
C1849 sky130_fd_sc_hd__nand2_8_4/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.05e-21
C1850 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# -4.66e-20
C1851 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# V_LOW -6.55e-19
C1852 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 0.00337f
C1853 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# V_GND 4.07e-19
C1854 sky130_fd_sc_hd__conb_1_25/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00207f
C1855 sky130_fd_sc_hd__conb_1_17/LO sky130_fd_sc_hd__conb_1_17/HI 0.00414f
C1856 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# -0.00139f
C1857 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# -2.32e-19
C1858 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 5.91e-20
C1859 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0034f
C1860 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 2.16e-20
C1861 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 1.58e-21
C1862 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 1.02e-19
C1863 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 4.12e-19
C1864 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# V_GND 1.15e-19
C1865 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# sky130_fd_sc_hd__conb_1_13/HI 1.83e-19
C1866 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# V_GND -0.00365f
C1867 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# -6.29e-19
C1868 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_557_413# -3.67e-20
C1869 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# V_LOW 1.38e-19
C1870 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__nand2_8_9/Y 4.06e-21
C1871 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# -0.0201f
C1872 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# -0.0078f
C1873 sky130_fd_sc_hd__dfbbn_1_26/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 9.46e-20
C1874 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# V_GND 0.00367f
C1875 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# V_GND 0.00249f
C1876 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/Q_N -9.56e-20
C1877 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_70/A 2.71e-19
C1878 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 2.8e-19
C1879 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 5.93e-21
C1880 sky130_fd_sc_hd__inv_1_65/Y V_GND 0.265f
C1881 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 2.49e-19
C1882 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0.00104f
C1883 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand3_1_2/B 0.045f
C1884 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_557_413# 5.03e-19
C1885 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00457f
C1886 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# V_GND 0.0035f
C1887 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_56/Y 1.3e-19
C1888 sky130_fd_sc_hd__nand3_1_2/a_109_47# V_GND 2.21e-19
C1889 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1_70/A 0.00988f
C1890 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# V_GND 0.00144f
C1891 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# V_LOW 1.38e-19
C1892 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.38e-20
C1893 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# V_LOW 3.56e-20
C1894 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI -9.23e-19
C1895 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 0.0194f
C1896 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# V_GND -0.0105f
C1897 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# V_LOW -9.15e-19
C1898 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.01e-20
C1899 sky130_fd_sc_hd__dfbbn_1_44/a_581_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.49e-19
C1900 sky130_fd_sc_hd__inv_16_1/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 2.67e-20
C1901 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.15e-19
C1902 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_16/HI 6.16e-20
C1903 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.07e-19
C1904 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# V_GND 0.00114f
C1905 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.57e-21
C1906 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_20/LO 5.04e-21
C1907 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_41/HI 3.31e-19
C1908 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 0.0112f
C1909 sky130_fd_sc_hd__inv_1_19/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00261f
C1910 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# -0.00184f
C1911 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__dfbbn_1_20/a_941_21# -7.6e-19
C1912 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# -0.00263f
C1913 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# Reset 0.00202f
C1914 sky130_fd_sc_hd__conb_1_29/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0512f
C1915 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_95/A 0.0844f
C1916 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# V_GND 8.12e-19
C1917 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_891_329# 0.00313f
C1918 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# V_GND 2.03e-19
C1919 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/Q_N 2.04e-20
C1920 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_891_329# -0.00159f
C1921 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# -0.00486f
C1922 sky130_fd_sc_hd__inv_1_3/Y V_SENSE 0.0661f
C1923 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# V_GND 1.08e-19
C1924 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0819f
C1925 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# V_LOW -0.00338f
C1926 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# V_GND -0.00531f
C1927 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 8.98e-19
C1928 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_12/HI 3.71e-20
C1929 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__nand3_1_2/Y 2.37e-20
C1930 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__inv_1_54/Y 4.59e-21
C1931 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 0.0238f
C1932 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00225f
C1933 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0.0086f
C1934 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 4.4e-20
C1935 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 4.4e-20
C1936 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0.0086f
C1937 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00135f
C1938 FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_50/Y 6.24e-20
C1939 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__conb_1_22/HI 6.44e-20
C1940 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/Q_N 0.0323f
C1941 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.00268f
C1942 sky130_fd_sc_hd__conb_1_51/LO V_GND -0.0057f
C1943 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# -0.00336f
C1944 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# -3.79e-20
C1945 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00134f
C1946 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0279f
C1947 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 1.75e-19
C1948 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.0229f
C1949 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF0.Q 0.051f
C1950 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/Q_N -9.56e-20
C1951 sky130_fd_sc_hd__inv_1_8/Y V_GND 0.0628f
C1952 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI 3.02e-19
C1953 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 4.12e-20
C1954 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# 2.1e-21
C1955 sky130_fd_sc_hd__inv_1_71/Y Reset 1.85e-19
C1956 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 0.011f
C1957 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# V_LOW 2.26e-20
C1958 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# V_GND 6.73e-19
C1959 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 4.24e-19
C1960 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_15/Y 5.93e-21
C1961 sky130_fd_sc_hd__inv_1_50/Y V_LOW 0.387f
C1962 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__inv_1_12/Y 7.4e-19
C1963 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_1_65/Y 2.55e-21
C1964 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 1.34e-20
C1965 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 7.38e-21
C1966 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 3.82e-20
C1967 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 2.73e-19
C1968 sky130_fd_sc_hd__conb_1_9/LO FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0469f
C1969 sky130_fd_sc_hd__inv_1_90/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0145f
C1970 sky130_fd_sc_hd__nand3_1_1/Y sky130_fd_sc_hd__inv_1_65/Y 0.0687f
C1971 sky130_fd_sc_hd__nor2_1_0/Y V_GND -3.79e-19
C1972 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# sky130_fd_sc_hd__inv_1_12/Y 2.65e-19
C1973 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.01e-21
C1974 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.47e-19
C1975 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 0.00178f
C1976 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# -1.64e-19
C1977 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 3.11e-21
C1978 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 0.00323f
C1979 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# sky130_fd_sc_hd__inv_1_9/Y 1.72e-20
C1980 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# V_LOW 0.0247f
C1981 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.5e-19
C1982 sky130_fd_sc_hd__dfbbn_1_34/Q_N V_GND -0.00753f
C1983 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI 0.00336f
C1984 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_28/HI 0.309f
C1985 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_80/A 0.0548f
C1986 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# V_GND 0.0018f
C1987 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# V_LOW -0.00387f
C1988 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# V_GND -0.00291f
C1989 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 1.08e-19
C1990 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 2.44e-20
C1991 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 4.21e-20
C1992 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 1.28e-20
C1993 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 9.16e-19
C1994 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0594f
C1995 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00429f
C1996 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_381_47# -0.00441f
C1997 sky130_fd_sc_hd__dfbbn_1_42/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00217f
C1998 sky130_fd_sc_hd__conb_1_50/LO V_LOW 0.0638f
C1999 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.0188f
C2000 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__conb_1_15/LO 9.95e-20
C2001 sky130_fd_sc_hd__dfbbn_1_29/Q_N V_GND -5.19e-19
C2002 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.43e-20
C2003 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__conb_1_44/HI 6.08e-21
C2004 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00574f
C2005 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# V_GND 0.01f
C2006 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__conb_1_45/HI 0.0283f
C2007 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00477f
C2008 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.45e-20
C2009 sky130_fd_sc_hd__dfbbn_1_46/a_557_413# V_GND 2.69e-19
C2010 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.65e-21
C2011 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 6.79e-20
C2012 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00431f
C2013 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__conb_1_41/HI 3.29e-20
C2014 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.0037f
C2015 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# V_GND 7.43e-19
C2016 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0196f
C2017 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/Q_N -9.56e-20
C2018 sky130_fd_sc_hd__nand2_8_9/a_27_47# Reset 4.5e-19
C2019 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_557_413# 5.03e-19
C2020 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -4.98e-19
C2021 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_473_413# -0.0103f
C2022 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# -9.32e-20
C2023 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_75/A 0.0215f
C2024 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 8.4e-21
C2025 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 6.66e-19
C2026 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 9.05e-19
C2027 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.003f
C2028 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 3.99e-20
C2029 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00225f
C2030 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__conb_1_8/HI 1.67e-19
C2031 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# Reset 4.39e-20
C2032 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# -3.46e-20
C2033 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 1.42e-32
C2034 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__inv_2_0/Y 1.78e-19
C2035 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_381_47# -2.53e-20
C2036 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_1_98/Y 0.00168f
C2037 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# V_GND -0.00948f
C2038 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__conb_1_51/HI 0.019f
C2039 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_891_329# -2.2e-20
C2040 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# -1.55e-19
C2041 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 0.0016f
C2042 sky130_fd_sc_hd__dfbbn_1_36/Q_N V_GND 6.85e-19
C2043 sky130_fd_sc_hd__inv_1_63/Y sky130_fd_sc_hd__inv_1_9/Y 0.00382f
C2044 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.03e-19
C2045 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 8.69e-19
C2046 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.006f
C2047 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 1.13e-19
C2048 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 0.0108f
C2049 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 9.7e-20
C2050 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 0.167f
C2051 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.0511f
C2052 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__inv_1_12/Y 0.00219f
C2053 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_891_329# -0.00159f
C2054 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# -0.00588f
C2055 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 3.69e-20
C2056 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 3.29e-19
C2057 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_791_47# 3.69e-20
C2058 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 3.29e-19
C2059 sky130_fd_sc_hd__dfbbn_1_20/Q_N V_LOW -0.00509f
C2060 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 6.73e-20
C2061 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_61/Y 0.0641f
C2062 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_381_47# -3.79e-20
C2063 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# -0.00336f
C2064 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# 1.67e-21
C2065 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# V_LOW -0.321f
C2066 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0305f
C2067 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# -0.0996f
C2068 sky130_fd_sc_hd__conb_1_39/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00178f
C2069 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__conb_1_44/HI 6.95e-21
C2070 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__conb_1_47/HI 1.09e-19
C2071 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__conb_1_49/HI 6.9e-21
C2072 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 1.91f
C2073 sky130_fd_sc_hd__inv_1_58/Y V_GND 0.104f
C2074 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.0798f
C2075 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.57e-20
C2076 sky130_fd_sc_hd__dfbbn_1_15/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 2.96e-19
C2077 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# V_LOW 0.0269f
C2078 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.0025f
C2079 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# V_GND 0.0226f
C2080 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_1_3/a_113_47# 5.93e-19
C2081 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 6.71e-21
C2082 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# sky130_fd_sc_hd__inv_1_49/Y 3.12e-19
C2083 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 0.0115f
C2084 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 8.28e-21
C2085 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 4.94e-20
C2086 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# V_LOW -0.00266f
C2087 sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.281f
C2088 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_0/Y 4.06e-21
C2089 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__conb_1_23/HI 9.13e-20
C2090 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# V_LOW 0.00856f
C2091 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 8.74e-20
C2092 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# V_GND -0.0455f
C2093 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_76/A 0.0922f
C2094 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_35/HI 5.49e-21
C2095 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__conb_1_32/HI 9.97e-19
C2096 sky130_fd_sc_hd__dfbbn_1_1/Q_N V_GND -7.63e-19
C2097 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# V_GND 0.00793f
C2098 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__conb_1_2/LO 3.89e-20
C2099 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# 5.04e-19
C2100 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0.0135f
C2101 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 8.42e-19
C2102 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0.00193f
C2103 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 8.42e-19
C2104 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 0.00193f
C2105 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0.0135f
C2106 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_15/Y 0.0047f
C2107 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# V_GND 0.00755f
C2108 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 6.63e-19
C2109 sky130_fd_sc_hd__inv_1_109/Y V_LOW 0.083f
C2110 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/Q_N 4.47e-19
C2111 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_791_47# 6.86e-21
C2112 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 7.5e-21
C2113 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0276f
C2114 sky130_fd_sc_hd__dfbbn_1_23/Q_N RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0114f
C2115 sky130_fd_sc_hd__conb_1_18/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00293f
C2116 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__inv_1_15/Y 0.00178f
C2117 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# -1.44e-20
C2118 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0018f
C2119 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 6.45e-19
C2120 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.26e-19
C2121 sky130_fd_sc_hd__inv_1_101/Y V_GND 0.00874f
C2122 sky130_fd_sc_hd__dfbbn_1_42/Q_N FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.15e-19
C2123 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_103/Y 0.0297f
C2124 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00134f
C2125 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 5.23e-19
C2126 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# V_GND 2.47e-19
C2127 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__inv_1_108/Y 0.00185f
C2128 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__conb_1_27/HI 3.07e-19
C2129 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# -0.00813f
C2130 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# V_LOW 3.56e-20
C2131 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_61/Y 0.00739f
C2132 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.21e-19
C2133 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 8.74e-21
C2134 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0.00451f
C2135 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0039f
C2136 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 4.21e-21
C2137 sky130_fd_sc_hd__inv_16_1/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.186f
C2138 sky130_fd_sc_hd__fill_4_73/VPB V_GND 0.459f
C2139 Reset sky130_fd_sc_hd__conb_1_2/HI 0.0103f
C2140 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 4.15e-20
C2141 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.0017f
C2142 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__conb_1_47/LO 8.81e-20
C2143 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 1.31e-22
C2144 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.03e-19
C2145 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# -6.8e-19
C2146 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/Q_N -4.78e-20
C2147 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00238f
C2148 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__conb_1_48/LO 7.5e-19
C2149 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_23/Y -0.0024f
C2150 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 1.38e-21
C2151 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__conb_1_5/HI 5.08e-19
C2152 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 3.74e-20
C2153 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.45e-20
C2154 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# -1.44e-20
C2155 sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__inv_1_99/Y 0.0789f
C2156 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_35/a_941_21# -5.45e-20
C2157 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# V_GND 2.04e-19
C2158 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__conb_1_34/HI 4.14e-19
C2159 sky130_fd_sc_hd__conb_1_45/HI V_LOW 0.099f
C2160 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# -3.46e-20
C2161 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 2.62e-19
C2162 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.26e-20
C2163 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 9.81e-21
C2164 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 1.07e-20
C2165 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 8.81e-20
C2166 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 3.18e-20
C2167 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 1.36e-20
C2168 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 5.82e-20
C2169 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 9.65e-21
C2170 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 5.74e-19
C2171 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.0036f
C2172 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 3.13e-21
C2173 sky130_fd_sc_hd__dfbbn_1_17/a_557_413# V_LOW 3.56e-20
C2174 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 6e-21
C2175 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# 0.00238f
C2176 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.11e-20
C2177 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.17e-20
C2178 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# sky130_fd_sc_hd__inv_1_12/Y 6.42e-19
C2179 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 1.29e-19
C2180 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 9.93e-21
C2181 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__conb_1_33/LO 1.71e-19
C2182 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# -1.42e-32
C2183 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# -0.00592f
C2184 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 7.32e-22
C2185 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_2/HI 5.07e-19
C2186 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0298f
C2187 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00237f
C2188 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_14/LO 0.00126f
C2189 FALLING_COUNTER.COUNT_SUB_DFF11.Q V_LOW 0.898f
C2190 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 5.62e-21
C2191 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 2.95e-21
C2192 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00174f
C2193 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 1.34e-19
C2194 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF15.Q 0.119f
C2195 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 0.0254f
C2196 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# V_LOW 4.33e-20
C2197 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_68/A 0.141f
C2198 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_6/LO 0.00716f
C2199 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_103/Y 0.0244f
C2200 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_17/HI 0.347f
C2201 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# V_LOW 2.26e-20
C2202 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# sky130_fd_sc_hd__inv_1_8/Y 3.75e-21
C2203 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# V_LOW 2.94e-20
C2204 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# V_GND 1.48e-19
C2205 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.22e-19
C2206 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.33e-20
C2207 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_49/LO 0.00109f
C2208 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# 0.00154f
C2209 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__inv_1_100/Y 2.49e-19
C2210 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 0.0101f
C2211 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00986f
C2212 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/Q_N 1.56e-19
C2213 sky130_fd_sc_hd__conb_1_5/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0507f
C2214 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/Q_N 3.91e-19
C2215 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_11/HI 2.77e-20
C2216 RISING_COUNTER.COUNT_SUB_DFF7.Q V_GND 1.49f
C2217 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_12/HI 0.0853f
C2218 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# V_GND 2.42e-19
C2219 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 1.29e-20
C2220 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 1.42e-20
C2221 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 1.85e-20
C2222 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__conb_1_13/LO 2.72e-20
C2223 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_17/Y 2.22e-20
C2224 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# V_GND 0.00192f
C2225 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.69e-20
C2226 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# -0.0122f
C2227 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -1.61e-19
C2228 sky130_fd_sc_hd__nand2_1_2/a_113_47# V_GND 8.29e-21
C2229 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# V_GND 0.00132f
C2230 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 3.98e-19
C2231 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 3.98e-19
C2232 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_193_47# 1.63e-19
C2233 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_97/A 0.00737f
C2234 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__inv_1_15/Y 4.86e-19
C2235 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_93/Y 0.00163f
C2236 RISING_COUNTER.COUNT_SUB_DFF6.Q V_LOW 1.44f
C2237 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_557_413# 8.17e-19
C2238 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__inv_1_16/Y 0.0112f
C2239 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 0.00224f
C2240 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.07e-19
C2241 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_40/HI 0.191f
C2242 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__inv_1_103/Y 0.00367f
C2243 sky130_fd_sc_hd__dfbbn_1_16/Q_N FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0264f
C2244 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# sky130_fd_sc_hd__inv_1_108/Y 5.8e-19
C2245 sky130_fd_sc_hd__inv_1_33/Y V_GND 0.0725f
C2246 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# -0.00107f
C2247 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# V_GND 0.00587f
C2248 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# 1.44e-20
C2249 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0479f
C2250 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# -0.00869f
C2251 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_40/a_193_47# 0.00453f
C2252 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 1.33e-20
C2253 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__inv_1_47/Y 0.00592f
C2254 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 0.00685f
C2255 sky130_fd_sc_hd__inv_1_39/A V_LOW 0.668f
C2256 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 7.37e-20
C2257 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_68/A 1.26e-19
C2258 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 1.18e-19
C2259 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# sky130_fd_sc_hd__conb_1_35/HI 5.79e-19
C2260 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_76/A 0.00225f
C2261 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_88/Y 0.00438f
C2262 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 5.04e-19
C2263 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.25e-19
C2264 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.23e-20
C2265 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.03e-20
C2266 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.88e-20
C2267 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_39/LO 1.15e-19
C2268 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.65e-21
C2269 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00194f
C2270 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.2e-20
C2271 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0403f
C2272 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__conb_1_0/HI 2.29e-19
C2273 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 5.44e-19
C2274 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__conb_1_5/HI 6.61e-20
C2275 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.77e-19
C2276 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.69e-19
C2277 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__inv_1_58/Y 1.75e-21
C2278 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 8.02e-20
C2279 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 5.88e-21
C2280 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# 4.27e-20
C2281 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 6.93e-22
C2282 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00119f
C2283 sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__nand2_8_9/Y 0.00914f
C2284 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 1.61e-19
C2285 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.34e-21
C2286 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 2.74e-20
C2287 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/Q_N 9.65e-21
C2288 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__conb_1_33/HI 5.85e-19
C2289 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__conb_1_2/HI 4.72e-19
C2290 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -2.36e-19
C2291 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# -0.00344f
C2292 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00618f
C2293 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__inv_1_103/Y 0.00568f
C2294 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 9.29e-19
C2295 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00216f
C2296 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_95/A 3.41e-19
C2297 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 1.09e-19
C2298 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0603f
C2299 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 2.3e-20
C2300 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 1.84e-20
C2301 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 1e-19
C2302 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.95e-20
C2303 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_581_47# 0.0011f
C2304 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# 0.00176f
C2305 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.03e-21
C2306 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 0.00554f
C2307 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 3.72e-19
C2308 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# V_LOW 0.0268f
C2309 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# V_LOW 7.12e-19
C2310 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# V_LOW 2.26e-20
C2311 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_86/Y 1.03e-19
C2312 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 4.73e-20
C2313 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__conb_1_11/LO 0.0682f
C2314 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# V_LOW 0.00613f
C2315 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 3.45e-19
C2316 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 3.37e-19
C2317 sky130_fd_sc_hd__inv_1_19/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 3.82e-19
C2318 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 0.00448f
C2319 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# 5.62e-19
C2320 FALLING_COUNTER.COUNT_SUB_DFF9.Q V_GND 1.1f
C2321 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_76/A 0.00133f
C2322 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# -3.06e-20
C2323 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# -0.00631f
C2324 sky130_fd_sc_hd__conb_1_7/LO V_GND -0.00465f
C2325 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0255f
C2326 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.128f
C2327 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# 2.12e-19
C2328 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__inv_1_58/Y 0.0023f
C2329 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# V_LOW 0.00758f
C2330 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__inv_16_1/Y 3.37e-19
C2331 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.11e-19
C2332 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_557_413# 1.85e-19
C2333 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# -2.57e-20
C2334 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 0.00137f
C2335 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_93/A 0.345f
C2336 sky130_fd_sc_hd__nor2_1_0/a_109_297# V_LOW 1.5e-19
C2337 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 7.97e-19
C2338 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/Q_N 7.97e-19
C2339 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_1_15/Y 3.2e-21
C2340 FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_106/Y 0.33f
C2341 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_16_1/Y 0.107f
C2342 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# V_LOW 0.0279f
C2343 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_108/Y 0.00282f
C2344 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__inv_1_50/Y 3.4e-20
C2345 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# V_GND -0.00537f
C2346 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# V_GND 2.12e-19
C2347 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# V_LOW 0.014f
C2348 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# -1.6e-19
C2349 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# -5.54e-21
C2350 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 0.0341f
C2351 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0117f
C2352 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# V_GND 0.0017f
C2353 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# V_GND 0.00373f
C2354 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_21/HI 0.201f
C2355 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# -1.44e-20
C2356 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# 0.00321f
C2357 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# V_GND 1.67e-19
C2358 sky130_fd_sc_hd__dfbbn_1_32/Q_N FALLING_COUNTER.COUNT_SUB_DFF3.Q 2.4e-19
C2359 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__inv_1_4/Y 7.07e-20
C2360 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_647_21# -0.00782f
C2361 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00534f
C2362 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 3.27e-19
C2363 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__nand3_1_2/Y 0.0023f
C2364 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_34/A 0.0443f
C2365 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_1/Y 1.6e-19
C2366 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 5.12e-21
C2367 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_647_21# -0.00797f
C2368 Reset sky130_fd_sc_hd__inv_2_0/Y 0.0187f
C2369 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 0.00327f
C2370 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__inv_1_57/Y 8.07e-20
C2371 sky130_fd_sc_hd__dfbbn_1_6/Q_N FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0195f
C2372 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_49/HI 0.0361f
C2373 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# V_GND 2.07e-19
C2374 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_1_15/Y 7.59e-21
C2375 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__inv_1_59/Y 0.0456f
C2376 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# V_GND 0.00766f
C2377 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0138f
C2378 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# sky130_fd_sc_hd__inv_16_2/Y 3.08e-20
C2379 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.54e-20
C2380 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.591f
C2381 sky130_fd_sc_hd__inv_1_85/A Reset 0.488f
C2382 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 2.32e-20
C2383 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 8.97e-19
C2384 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.34e-19
C2385 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# V_LOW -0.0199f
C2386 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# V_GND 0.0061f
C2387 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__inv_1_21/Y 4.82e-19
C2388 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 0.00581f
C2389 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 7.36e-19
C2390 FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_16_2/Y 0.262f
C2391 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00244f
C2392 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.92e-20
C2393 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# sky130_fd_sc_hd__conb_1_33/HI 0.00199f
C2394 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 8.7e-20
C2395 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_24/HI 3.36e-19
C2396 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# -2.57e-20
C2397 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.76e-20
C2398 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.192f
C2399 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_647_21# -0.00122f
C2400 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# -0.00339f
C2401 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00624f
C2402 sky130_fd_sc_hd__conb_1_3/HI V_GND 0.044f
C2403 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00315f
C2404 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__inv_1_20/Y 2.78e-19
C2405 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_97/A 0.154f
C2406 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__conb_1_27/LO 4.69e-19
C2407 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__inv_1_62/Y 9.4e-19
C2408 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# -0.00133f
C2409 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# -0.00512f
C2410 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# V_GND 2.48e-19
C2411 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.01e-21
C2412 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 1.93e-19
C2413 sky130_fd_sc_hd__inv_1_10/Y sky130_fd_sc_hd__conb_1_0/HI 0.037f
C2414 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.00122f
C2415 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00736f
C2416 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.96e-20
C2417 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# 5.32e-19
C2418 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__inv_1_17/Y 2.44e-19
C2419 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# V_LOW 0.0174f
C2420 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.39e-19
C2421 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 2.96e-20
C2422 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 8.02e-20
C2423 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 3.55e-19
C2424 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__conb_1_38/LO 0.0144f
C2425 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.00515f
C2426 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.67e-19
C2427 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0687f
C2428 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__nand3_1_1/a_193_47# 6.99e-19
C2429 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# V_LOW -0.00103f
C2430 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_21/HI 0.13f
C2431 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# V_LOW -2.57e-19
C2432 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 9.18e-19
C2433 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__inv_1_108/Y 9.89e-22
C2434 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.031f
C2435 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_16_2/Y 0.00749f
C2436 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_0/Y 0.33f
C2437 sky130_fd_sc_hd__inv_1_70/Y Reset 7.53e-19
C2438 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.248f
C2439 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# V_LOW 0.00496f
C2440 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# V_GND -0.0051f
C2441 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_105/Y 1.19e-20
C2442 FALLING_COUNTER.COUNT_SUB_DFF8.Q V_LOW 2.54f
C2443 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# -9.32e-20
C2444 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0196f
C2445 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0128f
C2446 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# V_GND 0.0019f
C2447 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_21/HI 2.29e-19
C2448 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF1.Q 2.12e-19
C2449 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/Q_N 0.0036f
C2450 RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_24/HI 0.00218f
C2451 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# V_LOW 2.26e-20
C2452 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# V_GND 0.00481f
C2453 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_581_47# -2.6e-20
C2454 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# CLOCK_GEN.SR_Op.Q 1.36e-19
C2455 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0.00133f
C2456 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.037f
C2457 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 3.11e-19
C2458 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 1.86e-20
C2459 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__conb_1_46/HI 1.7e-20
C2460 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00992f
C2461 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_581_47# -2.6e-20
C2462 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.45e-19
C2463 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.0449f
C2464 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.69e-20
C2465 sky130_fd_sc_hd__conb_1_36/LO FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0588f
C2466 sky130_fd_sc_hd__inv_1_61/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0453f
C2467 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__conb_1_49/HI 4.59e-19
C2468 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00109f
C2469 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0514f
C2470 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__inv_1_15/Y 1.6e-19
C2471 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00175f
C2472 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# V_GND 0.00629f
C2473 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 1.77e-20
C2474 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__inv_1_112/Y 0.00265f
C2475 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 1.89e-19
C2476 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.0099f
C2477 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00258f
C2478 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF14.Q 0.427f
C2479 sky130_fd_sc_hd__inv_16_2/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.324f
C2480 sky130_fd_sc_hd__dfbbn_1_28/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 3.01e-20
C2481 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 0.00415f
C2482 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_557_413# 2.55e-19
C2483 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_0/Q_N 5.11e-19
C2484 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.11f
C2485 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# -0.00827f
C2486 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -0.00117f
C2487 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -9.88e-20
C2488 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# V_LOW -0.00604f
C2489 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# V_GND 0.00173f
C2490 sky130_fd_sc_hd__conb_1_47/LO FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0101f
C2491 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_891_329# -2.2e-20
C2492 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# -4.1e-19
C2493 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 1.55e-20
C2494 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__conb_1_30/HI 0.00126f
C2495 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 0.00144f
C2496 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_5/Y 0.562f
C2497 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_96/Y 0.00342f
C2498 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0136f
C2499 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# -0.0489f
C2500 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00284f
C2501 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# -0.00138f
C2502 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.00193f
C2503 sky130_fd_sc_hd__dfbbn_1_41/Q_N RISING_COUNTER.COUNT_SUB_DFF2.Q 7.06e-21
C2504 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.46e-19
C2505 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 6.31e-19
C2506 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 0.0237f
C2507 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_12/Q_N 7.97e-21
C2508 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# -2.56e-19
C2509 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# -2.37e-19
C2510 sky130_fd_sc_hd__conb_1_20/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 6.54e-20
C2511 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.71e-19
C2512 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# -0.00832f
C2513 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -9.88e-20
C2514 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# -0.00125f
C2515 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 6.5e-20
C2516 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0319f
C2517 sky130_fd_sc_hd__dfbbn_1_48/Q_N RISING_COUNTER.COUNT_SUB_DFF6.Q 4.87e-20
C2518 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_94/A 0.291f
C2519 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0517f
C2520 FULL_COUNTER.COUNT_SUB_DFF8.Q V_GND 3.21f
C2521 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# sky130_fd_sc_hd__inv_1_17/Y 7.36e-20
C2522 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 0.00154f
C2523 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 5.85e-21
C2524 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# V_LOW -0.00363f
C2525 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_381_47# -0.00538f
C2526 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# -6.22e-19
C2527 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# -0.00117f
C2528 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.56e-19
C2529 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 8.31e-20
C2530 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.92e-19
C2531 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 4.05e-19
C2532 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__inv_1_11/Y 2.57e-20
C2533 CLOCK_GEN.SR_Op.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 1.03f
C2534 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_63/Y 0.244f
C2535 sky130_fd_sc_hd__dfbbn_1_39/a_581_47# sky130_fd_sc_hd__inv_1_108/Y 2.32e-20
C2536 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_1_5/Y 1.07e-21
C2537 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00762f
C2538 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 6.57e-22
C2539 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 4.14e-20
C2540 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_1_90/Y 0.00373f
C2541 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.04e-19
C2542 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__inv_1_9/Y 0.00837f
C2543 sky130_fd_sc_hd__dfbbn_1_26/Q_N V_GND -0.00726f
C2544 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__conb_1_9/LO 3.43e-20
C2545 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__inv_1_11/Y 0.0114f
C2546 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/Q_N -4.78e-20
C2547 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/Q_N 0.0253f
C2548 sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00278f
C2549 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# V_GND 8.4e-19
C2550 sky130_fd_sc_hd__dfbbn_1_31/Q_N V_GND -0.00169f
C2551 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 1.63e-19
C2552 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# V_LOW 0.0012f
C2553 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_891_329# -2.2e-20
C2554 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -0.00915f
C2555 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI 7.25e-22
C2556 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__conb_1_37/HI -0.002f
C2557 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.48e-19
C2558 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# V_GND 0.00174f
C2559 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_6/HI 3.23e-19
C2560 FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_12/Y 0.171f
C2561 FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_20/Y 1.16e-20
C2562 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 0.0012f
C2563 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 0.0402f
C2564 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 1.21e-19
C2565 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0.0498f
C2566 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 4.55e-20
C2567 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0158f
C2568 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 5.44e-19
C2569 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 3.65e-21
C2570 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 6.11e-21
C2571 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 1.64e-20
C2572 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.36e-19
C2573 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_381_47# -3.05e-20
C2574 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# -0.00336f
C2575 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 5.71e-19
C2576 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.15e-21
C2577 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__nand2_8_2/A 4.66e-19
C2578 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_1_15/Y 4.38e-19
C2579 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_1_19/Y 1.56e-20
C2580 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 2.62e-19
C2581 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_37/LO 0.00289f
C2582 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 2.76e-20
C2583 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 8.79e-22
C2584 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 2.21e-19
C2585 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 6.46e-19
C2586 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# V_GND 0.00202f
C2587 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0264f
C2588 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_12/HI 0.442f
C2589 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# -0.00385f
C2590 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# -1.42e-32
C2591 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__conb_1_40/HI 1.09e-19
C2592 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_85/Y 0.135f
C2593 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 8.86e-21
C2594 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 9.95e-21
C2595 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# 8.86e-21
C2596 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# 9.95e-21
C2597 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_37/HI 0.00528f
C2598 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 7.88e-20
C2599 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_6/HI 3.57e-21
C2600 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.19e-20
C2601 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 8.86e-21
C2602 sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__inv_2_0/Y 0.00178f
C2603 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 4.5e-20
C2604 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_46/HI 0.011f
C2605 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nand3_1_2/B 5.52e-19
C2606 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 1.11e-20
C2607 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0294f
C2608 sky130_fd_sc_hd__inv_1_55/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0485f
C2609 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_41/LO 1.49e-19
C2610 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_1_59/Y 1.76e-19
C2611 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 9.48e-19
C2612 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_791_47# 9.26e-20
C2613 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 3.77e-21
C2614 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.00138f
C2615 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 9.2e-20
C2616 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.98e-19
C2617 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00545f
C2618 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00378f
C2619 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -1.66e-19
C2620 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/Q_N -9.56e-20
C2621 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.59e-19
C2622 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_51/LO 0.00154f
C2623 CLOCK_GEN.SR_Op.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0289f
C2624 RISING_COUNTER.COUNT_SUB_DFF2.Q Reset 1.98e-19
C2625 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.75e-20
C2626 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_1_99/Y 8.47e-19
C2627 sky130_fd_sc_hd__inv_1_97/A V_LOW 0.188f
C2628 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 5.18e-19
C2629 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# V_LOW -0.00212f
C2630 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1_23/LO 0.00158f
C2631 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.182f
C2632 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 3.95e-19
C2633 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# 5.83e-19
C2634 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.86e-19
C2635 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 4.06e-21
C2636 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 1.55e-20
C2637 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__conb_1_8/HI 0.0132f
C2638 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__conb_1_6/HI 0.00214f
C2639 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_5/HI 0.0382f
C2640 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__nand3_1_0/Y 4.11e-20
C2641 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 1.67e-20
C2642 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# sky130_fd_sc_hd__inv_1_11/Y 4.29e-20
C2643 FALLING_COUNTER.COUNT_SUB_DFF13.Q V_LOW 2.67f
C2644 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 0.00421f
C2645 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 3.77e-19
C2646 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# CLOCK_GEN.SR_Op.Q 8.73e-20
C2647 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__inv_1_62/Y 0.00186f
C2648 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0111f
C2649 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_68/A 0.0661f
C2650 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# V_LOW -0.0136f
C2651 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# CLOCK_GEN.SR_Op.Q 0.0342f
C2652 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 0.00344f
C2653 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00344f
C2654 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 7.7e-21
C2655 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.63e-21
C2656 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_47/Y 0.00194f
C2657 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# sky130_fd_sc_hd__inv_1_90/Y 1.07e-21
C2658 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 9.09e-19
C2659 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_1_16/Y 0.0208f
C2660 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_64/A 0.13f
C2661 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.421f
C2662 sky130_fd_sc_hd__dfbbn_1_39/a_557_413# V_GND 1.9e-19
C2663 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__conb_1_6/HI 1.85e-21
C2664 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00292f
C2665 sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 3.37e-19
C2666 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 1.36e-19
C2667 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0141f
C2668 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# -1.42e-32
C2669 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# -0.00592f
C2670 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__conb_1_31/HI 0.00311f
C2671 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__conb_1_31/HI 4.03e-21
C2672 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 5.9e-19
C2673 sky130_fd_sc_hd__inv_1_18/Y V_LOW 0.998f
C2674 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__conb_1_37/HI -4.01e-20
C2675 sky130_fd_sc_hd__dfbbn_1_19/Q_N V_GND -8.3e-19
C2676 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 1.67e-19
C2677 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 5.41e-19
C2678 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.325f
C2679 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 0.00248f
C2680 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__conb_1_13/HI 0.0291f
C2681 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_14/LO 0.012f
C2682 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 8.52e-21
C2683 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# V_GND 0.00972f
C2684 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 0.0015f
C2685 sky130_fd_sc_hd__nand2_8_3/A V_LOW 0.175f
C2686 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_66/Y 3.71e-20
C2687 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_1_108/Y 4.43e-21
C2688 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 0.0019f
C2689 FULL_COUNTER.COUNT_SUB_DFF0.Q V_GND 1.26f
C2690 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_42/HI 0.00991f
C2691 sky130_fd_sc_hd__inv_1_40/A sky130_fd_sc_hd__inv_1_43/A 0.00133f
C2692 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/Q_N 2.12e-19
C2693 sky130_fd_sc_hd__dfbbn_1_46/Q_N FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0145f
C2694 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__conb_1_27/HI 3.93e-20
C2695 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_791_47# 2.38e-20
C2696 sky130_fd_sc_hd__inv_1_81/Y V_GND 0.0851f
C2697 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/Q_N -1.39e-35
C2698 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.1e-19
C2699 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# sky130_fd_sc_hd__conb_1_40/HI 5.9e-19
C2700 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__inv_16_1/Y 8.09e-19
C2701 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_21/HI 0.0189f
C2702 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# 1.52e-19
C2703 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0.00295f
C2704 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_57/Y 0.159f
C2705 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_26/HI 0.00116f
C2706 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__conb_1_34/LO 0.0144f
C2707 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__inv_1_58/Y 1.63e-20
C2708 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.11e-20
C2709 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_1_9/Y 4.79e-20
C2710 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.155f
C2711 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_23/HI 0.0311f
C2712 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/Q_N -9.56e-20
C2713 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 4.21e-21
C2714 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 3.36e-20
C2715 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# V_LOW 0.00794f
C2716 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 9.36e-20
C2717 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__conb_1_12/HI 3.66e-19
C2718 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 0.00483f
C2719 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.7e-22
C2720 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_25/HI -7.19e-19
C2721 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/Q_N -9.56e-20
C2722 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00102f
C2723 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.05e-20
C2724 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 5.53e-20
C2725 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 6.09e-20
C2726 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# 2.25e-19
C2727 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 6.12e-20
C2728 sky130_fd_sc_hd__inv_1_93/A RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00529f
C2729 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 5.73e-19
C2730 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 0.00104f
C2731 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 7.48e-20
C2732 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# -0.0127f
C2733 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__inv_1_62/Y 1.16e-19
C2734 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_7/Y 2.6e-20
C2735 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# V_LOW -6.55e-19
C2736 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# CLOCK_GEN.SR_Op.Q 0.00144f
C2737 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 7.34e-19
C2738 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_581_47# 1.08e-20
C2739 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 3.8e-19
C2740 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__conb_1_12/HI 1.26e-19
C2741 sky130_fd_sc_hd__inv_1_109/Y FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00403f
C2742 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 3.94e-21
C2743 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 7.38e-21
C2744 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_791_47# 3.16e-19
C2745 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__inv_1_16/Y 0.0324f
C2746 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_93/A 7.56e-21
C2747 sky130_fd_sc_hd__conb_1_16/HI V_LOW 0.0274f
C2748 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__inv_1_54/Y 1.07e-20
C2749 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_76/A 0.042f
C2750 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 2.53e-19
C2751 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.63e-20
C2752 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 3.88e-19
C2753 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00334f
C2754 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.00401f
C2755 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 9.08e-19
C2756 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 3.22e-19
C2757 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.14e-19
C2758 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# V_LOW 0.0134f
C2759 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__conb_1_26/HI 3.65e-19
C2760 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0548f
C2761 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 7.19e-21
C2762 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# 2.51e-22
C2763 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__inv_1_72/A 0.0434f
C2764 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__nand3_1_1/Y 4.44e-19
C2765 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__inv_1_18/Y 0.0209f
C2766 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 1.06e-21
C2767 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__conb_1_6/HI -5.28e-19
C2768 sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# V_GND 8.05e-19
C2769 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# 4.24e-21
C2770 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_75/A 4.43e-21
C2771 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00224f
C2772 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 0.0126f
C2773 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 7.24e-19
C2774 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__inv_1_19/Y 1.96e-21
C2775 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# CLOCK_GEN.SR_Op.Q 3.99e-20
C2776 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__conb_1_42/HI 9.86e-19
C2777 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__conb_1_22/HI 4.28e-20
C2778 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# V_LOW 0.0186f
C2779 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_45/HI 3.23e-20
C2780 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# 0.00306f
C2781 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# V_GND 0.00461f
C2782 FULL_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0218f
C2783 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.05e-19
C2784 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00109f
C2785 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 5.18e-21
C2786 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF3.Q 2.55e-20
C2787 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.57e-20
C2788 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# sky130_fd_sc_hd__conb_1_21/HI 5.34e-19
C2789 sky130_fd_sc_hd__conb_1_9/LO V_LOW 0.093f
C2790 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00996f
C2791 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.00122f
C2792 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 1.34e-19
C2793 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_119/Y 0.00813f
C2794 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_50/a_941_21# 9.41e-22
C2795 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_38/LO 1.08e-19
C2796 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# -4.37e-20
C2797 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# -0.00216f
C2798 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# -6.22e-19
C2799 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 8.36e-19
C2800 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# -4.66e-20
C2801 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 7.72e-21
C2802 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_1_6/Y 0.00378f
C2803 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.00391f
C2804 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 7.31e-21
C2805 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00596f
C2806 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_18/HI 0.00242f
C2807 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_8_7/a_27_47# 2.99e-19
C2808 sky130_fd_sc_hd__inv_1_119/Y sky130_fd_sc_hd__nand2_1_0/Y 0.0284f
C2809 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# sky130_fd_sc_hd__inv_1_98/Y 3.21e-19
C2810 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# V_GND -0.0089f
C2811 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__conb_1_18/HI 0.0369f
C2812 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# V_GND 0.00484f
C2813 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_23/HI 3.21e-19
C2814 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__conb_1_23/HI 0.0618f
C2815 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# V_GND 0.00583f
C2816 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_791_47# 4.95e-20
C2817 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 6.64e-20
C2818 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 0.0086f
C2819 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.92f
C2820 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 1.31e-20
C2821 sky130_fd_sc_hd__inv_1_95/Y Reset 0.0032f
C2822 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__conb_1_12/HI 6.22e-19
C2823 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 9.81e-19
C2824 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 0.00232f
C2825 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__conb_1_25/HI -2.07e-19
C2826 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__inv_1_106/Y 5.15e-19
C2827 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_473_413# -3.86e-20
C2828 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_941_21# -1.03e-19
C2829 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__conb_1_16/HI 0.00561f
C2830 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# 0.00406f
C2831 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.007f
C2832 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__nand3_1_2/B 3.96e-20
C2833 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_12/HI 0.00133f
C2834 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 1.58e-20
C2835 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 1.46e-20
C2836 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand3_1_2/B 1.08e-20
C2837 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 0.0906f
C2838 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 2.16e-20
C2839 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 4.3e-21
C2840 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 4.97e-19
C2841 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__conb_1_22/HI 4.07e-19
C2842 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_97/Y 2.06e-19
C2843 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# -0.0185f
C2844 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -6.4e-19
C2845 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0218f
C2846 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_41/a_941_21# 2.93e-20
C2847 sky130_fd_sc_hd__conb_1_21/HI V_LOW 0.108f
C2848 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__conb_1_16/HI 0.001f
C2849 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__inv_1_18/Y 1.59e-20
C2850 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.85e-19
C2851 sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# V_LOW 2.94e-20
C2852 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.75e-19
C2853 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_5/Y 0.0255f
C2854 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# V_LOW 0.0261f
C2855 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_12/HI 0.00232f
C2856 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0459f
C2857 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 7.55e-20
C2858 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.12e-20
C2859 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# V_LOW -0.00371f
C2860 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.55e-19
C2861 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# -4.66e-20
C2862 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# -3.79e-20
C2863 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__conb_1_6/HI 0.00218f
C2864 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# V_GND 0.015f
C2865 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0112f
C2866 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 0.0069f
C2867 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 6.9e-20
C2868 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00274f
C2869 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_76/A 1.82e-20
C2870 sky130_fd_sc_hd__inv_1_100/Y sky130_fd_sc_hd__inv_1_101/Y 0.0334f
C2871 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# 1.67e-21
C2872 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__nand2_8_9/Y 4.36e-19
C2873 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1_22/HI 0.0373f
C2874 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# CLOCK_GEN.SR_Op.Q 5.24e-19
C2875 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.3e-19
C2876 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_18/Y 0.581f
C2877 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__conb_1_12/LO 0.00189f
C2878 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 0.00798f
C2879 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# -3.86e-20
C2880 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# -3.07e-19
C2881 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# V_LOW 5.15e-20
C2882 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__inv_1_57/Y 7.37e-19
C2883 sky130_fd_sc_hd__conb_1_17/HI V_GND 0.822f
C2884 sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# V_GND 6.67e-19
C2885 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.7e-19
C2886 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__inv_1_99/Y 2.55e-21
C2887 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0116f
C2888 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# V_GND 2.35e-19
C2889 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# V_LOW 4.8e-20
C2890 sky130_fd_sc_hd__inv_1_56/Y RISING_COUNTER.COUNT_SUB_DFF2.Q 2.53e-19
C2891 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0388f
C2892 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 7.73e-19
C2893 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# V_LOW 4.8e-20
C2894 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__conb_1_35/HI 0.0113f
C2895 sky130_fd_sc_hd__conb_1_46/HI V_LOW 0.045f
C2896 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# V_GND 4.99e-19
C2897 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__inv_16_0/Y 4.59e-19
C2898 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 5.77e-20
C2899 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF14.Q 6.06e-19
C2900 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 0.00104f
C2901 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.17e-20
C2902 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 4.34e-20
C2903 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_10/Y 0.0503f
C2904 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 7.05e-19
C2905 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 1.03e-19
C2906 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 4.69e-19
C2907 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 3.57e-20
C2908 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__conb_1_40/HI 9.4e-19
C2909 sky130_fd_sc_hd__inv_2_0/A V_SENSE 3.32e-19
C2910 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00408f
C2911 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0399f
C2912 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 0.00256f
C2913 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_1_103/Y 0.00923f
C2914 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_41/LO 0.012f
C2915 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__conb_1_44/HI 4.39e-19
C2916 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.89e-21
C2917 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.81e-19
C2918 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# V_GND 3.39e-19
C2919 sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 0.449f
C2920 sky130_fd_sc_hd__conb_1_32/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.127f
C2921 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__nand3_1_0/Y 3.94e-19
C2922 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__conb_1_18/HI 0.0313f
C2923 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0.00492f
C2924 sky130_fd_sc_hd__dfbbn_1_38/a_581_47# V_GND 2.58e-19
C2925 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__conb_1_38/HI 0.00502f
C2926 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# V_LOW 1.38e-19
C2927 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_51/LO 0.0501f
C2928 sky130_fd_sc_hd__dfbbn_1_50/a_581_47# V_GND 2.87e-19
C2929 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0.00106f
C2930 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# V_LOW -0.00389f
C2931 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_1_23/Y 1.91e-19
C2932 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 1.41e-19
C2933 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# 7.82e-20
C2934 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 1.2e-19
C2935 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# sky130_fd_sc_hd__conb_1_28/HI -0.0123f
C2936 sky130_fd_sc_hd__inv_2_0/Y V_HIGH 1.54f
C2937 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/Q_N 0.00255f
C2938 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_9/LO 4.65e-19
C2939 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0393f
C2940 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# -2.57e-20
C2941 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# -3.79e-20
C2942 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# -0.00336f
C2943 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_94/A 0.048f
C2944 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_37/HI 0.00268f
C2945 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__conb_1_21/HI 6.32e-20
C2946 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__conb_1_12/HI 9.04e-19
C2947 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.73e-19
C2948 sky130_fd_sc_hd__inv_1_75/Y V_GND 0.0578f
C2949 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_97/Y 4.75e-20
C2950 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_381_47# -3.79e-20
C2951 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# -4.66e-20
C2952 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__conb_1_51/HI 1.12e-19
C2953 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# V_LOW -0.00121f
C2954 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 0.0254f
C2955 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# V_GND 9.25e-19
C2956 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.69f
C2957 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__conb_1_22/HI 2.43e-19
C2958 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# V_GND 7.5e-19
C2959 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# -6.8e-19
C2960 sky130_fd_sc_hd__nand2_8_6/a_27_47# V_LOW -0.00697f
C2961 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_1_54/Y 5.85e-22
C2962 Reset FULL_COUNTER.COUNT_SUB_DFF1.Q 2.68e-19
C2963 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__conb_1_16/HI -2.07e-19
C2964 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.0159f
C2965 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# V_LOW 0.0171f
C2966 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# -3.86e-20
C2967 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# -0.00442f
C2968 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 0.00561f
C2969 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 0.0134f
C2970 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_40/HI 0.00205f
C2971 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 3.82e-21
C2972 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# sky130_fd_sc_hd__inv_1_102/Y 4.15e-20
C2973 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.09e-20
C2974 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.46e-20
C2975 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__conb_1_6/HI -2.17e-19
C2976 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# V_GND -0.0036f
C2977 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0291f
C2978 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 1.45e-19
C2979 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00243f
C2980 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 1.41e-20
C2981 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 2.58e-20
C2982 sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__nand2_8_9/Y 0.0896f
C2983 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__inv_16_2/Y 0.0167f
C2984 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 3.08e-20
C2985 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 2.73e-20
C2986 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00287f
C2987 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__conb_1_12/LO 0.00251f
C2988 sky130_fd_sc_hd__inv_1_110/Y V_LOW 0.0816f
C2989 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# -2.57e-20
C2990 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__conb_1_18/HI 3.85e-19
C2991 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# V_GND 0.00956f
C2992 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00358f
C2993 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_557_413# -3.67e-20
C2994 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# -0.00717f
C2995 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_891_329# -2.46e-19
C2996 sky130_fd_sc_hd__dfbbn_1_45/Q_N FALLING_COUNTER.COUNT_SUB_DFF7.Q 2.19e-20
C2997 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0496f
C2998 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.73e-19
C2999 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 0.00528f
C3000 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.131f
C3001 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# V_LOW 0.00666f
C3002 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# -0.00199f
C3003 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# -0.00527f
C3004 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# Reset 2.22e-19
C3005 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 5.16e-19
C3006 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__conb_1_40/HI -2.65e-20
C3007 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0084f
C3008 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00482f
C3009 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 5.93e-19
C3010 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/Q_N -9.56e-20
C3011 RISING_COUNTER.COUNT_SUB_DFF0.Q V_GND 5.84f
C3012 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__nand3_1_0/Y 4.85e-21
C3013 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.34e-19
C3014 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_1_58/Y 0.00289f
C3015 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# -0.0496f
C3016 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__conb_1_35/HI 6.84e-21
C3017 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0222f
C3018 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 1.33e-19
C3019 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__conb_1_38/HI 8.57e-19
C3020 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_97/Y 0.356f
C3021 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_76/A 0.0415f
C3022 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# V_GND 0.0174f
C3023 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_53/Y 5.1e-20
C3024 sky130_fd_sc_hd__conb_1_5/LO V_LOW 0.0964f
C3025 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__conb_1_11/LO 1.38e-21
C3026 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_12/LO 3.73e-21
C3027 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 7.37e-19
C3028 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.34e-19
C3029 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_791_47# 2.47e-19
C3030 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__inv_16_0/Y 0.00696f
C3031 sky130_fd_sc_hd__conb_1_11/HI V_LOW 0.125f
C3032 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/Q_N 8.96e-21
C3033 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_74/Y 0.0146f
C3034 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_1_7/Y 1.26e-19
C3035 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_13/HI 6.45e-19
C3036 sky130_fd_sc_hd__conb_1_11/HI sky130_fd_sc_hd__conb_1_13/HI 4.03e-21
C3037 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_47/Y 2.65e-20
C3038 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF4.Q 8.27e-21
C3039 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_37/HI 0.00156f
C3040 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_85/Y 2.26e-19
C3041 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 2.48e-20
C3042 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 2.19e-19
C3043 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 1.22e-19
C3044 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__conb_1_12/HI 0.00987f
C3045 CLOCK_GEN.SR_Op.Q V_LOW 7.59f
C3046 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.47e-19
C3047 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_37/LO 0.00348f
C3048 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# -0.0197f
C3049 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_891_329# -2.46e-19
C3050 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_557_413# -3.67e-20
C3051 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__inv_1_57/Y 0.00348f
C3052 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__nand3_1_2/B 0.0319f
C3053 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 5.6e-21
C3054 sky130_fd_sc_hd__nand2_8_3/a_27_47# V_GND -3.26e-19
C3055 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__conb_1_22/HI 4.38e-20
C3056 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 0.00136f
C3057 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__conb_1_48/HI 2.17e-19
C3058 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_55/Y 4.59e-19
C3059 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0271f
C3060 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 0.00205f
C3061 sky130_fd_sc_hd__nand2_8_8/a_27_47# V_LOW -0.0116f
C3062 Reset sky130_fd_sc_hd__inv_1_72/A 0.0481f
C3063 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# V_LOW -0.0038f
C3064 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# V_LOW 2.26e-20
C3065 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 3.7e-19
C3066 sky130_fd_sc_hd__inv_1_75/A V_LOW 0.841f
C3067 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 1.44e-19
C3068 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 6.4e-20
C3069 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 1.81e-19
C3070 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# -8.41e-19
C3071 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 0.00396f
C3072 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__inv_1_57/Y 0.0452f
C3073 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__nand3_1_1/Y 6.25e-21
C3074 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.109f
C3075 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 8.29e-19
C3076 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.86e-19
C3077 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 2.39e-19
C3078 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.24e-20
C3079 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 1.86e-19
C3080 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 2.39e-19
C3081 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.24e-20
C3082 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_101/Y -3.93e-24
C3083 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00161f
C3084 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00842f
C3085 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0133f
C3086 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/Q_N 9.65e-21
C3087 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 3.73e-20
C3088 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__inv_1_93/A 0.0022f
C3089 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.127f
C3090 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 0.0016f
C3091 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_1_55/Y 3.32e-20
C3092 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_28/Y 1.6e-20
C3093 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 8.86e-19
C3094 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 5.69e-19
C3095 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__nand3_1_1/Y 8.41e-20
C3096 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 0.0353f
C3097 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# V_GND 5.57e-19
C3098 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# V_GND 0.00215f
C3099 sky130_fd_sc_hd__dfbbn_1_50/Q_N FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0352f
C3100 sky130_fd_sc_hd__dfbbn_1_0/Q_N FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0193f
C3101 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__conb_1_32/HI -1.32e-19
C3102 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# V_LOW 2.26e-20
C3103 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_647_21# 0.00486f
C3104 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__conb_1_9/LO 0.00139f
C3105 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0197f
C3106 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__nand3_1_2/Y 0.00987f
C3107 sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__inv_1_71/Y 3.52e-19
C3108 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__conb_1_0/HI 0.0199f
C3109 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# V_GND -0.155f
C3110 sky130_fd_sc_hd__fill_4_85/VPB V_GND 0.422f
C3111 sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__inv_1_80/A 2.11e-19
C3112 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# sky130_fd_sc_hd__inv_1_58/Y 5.8e-19
C3113 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_61/Y 0.0236f
C3114 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# V_GND -0.00447f
C3115 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_66/Y 5.57e-20
C3116 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# CLOCK_GEN.SR_Op.Q 8.11e-21
C3117 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__conb_1_34/HI 0.0174f
C3118 sky130_fd_sc_hd__conb_1_45/LO sky130_fd_sc_hd__conb_1_45/HI 0.00126f
C3119 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__nand2_8_3/Y 0.00633f
C3120 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0247f
C3121 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.049f
C3122 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.28e-20
C3123 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# -9.32e-20
C3124 sky130_fd_sc_hd__inv_1_71/A V_GND 1.01f
C3125 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 7.28e-21
C3126 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_381_47# -0.00375f
C3127 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# 1.6e-21
C3128 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 5.15e-21
C3129 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 1.02e-19
C3130 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.52e-19
C3131 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0577f
C3132 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0067f
C3133 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__conb_1_9/HI 0.00246f
C3134 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.51e-19
C3135 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_63/Y 0.0167f
C3136 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_45/HI 0.273f
C3137 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_22/HI 0.0184f
C3138 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 2.84e-19
C3139 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_581_47# 4.99e-19
C3140 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# sky130_fd_sc_hd__conb_1_48/HI 6.48e-20
C3141 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__conb_1_5/LO 2.51e-20
C3142 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 8.17e-19
C3143 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00385f
C3144 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# -0.00336f
C3145 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# V_LOW -0.00389f
C3146 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0413f
C3147 sky130_fd_sc_hd__conb_1_43/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0261f
C3148 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_80/A 0.0156f
C3149 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# 4.18e-19
C3150 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 7.41e-19
C3151 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/Q_N 0.00762f
C3152 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_1_22/Y 1.78e-21
C3153 sky130_fd_sc_hd__conb_1_42/HI V_GND -0.111f
C3154 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_1_60/Y 0.00947f
C3155 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 8.82e-21
C3156 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 2.07e-21
C3157 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 2.42e-20
C3158 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_791_47# 2.42e-20
C3159 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 2.07e-21
C3160 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 8.82e-21
C3161 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_40/LO 8.84e-20
C3162 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__conb_1_5/HI 0.00137f
C3163 sky130_fd_sc_hd__conb_1_34/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 5.27e-19
C3164 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.08e-20
C3165 sky130_fd_sc_hd__inv_1_90/Y sky130_fd_sc_hd__inv_1_59/Y 0.00258f
C3166 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0144f
C3167 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 1.75e-19
C3168 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.00121f
C3169 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 5.12e-20
C3170 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00177f
C3171 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 0.126f
C3172 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# V_LOW 0.0025f
C3173 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 5.87e-20
C3174 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__inv_1_71/Y 0.00157f
C3175 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# V_LOW 3.56e-20
C3176 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0345f
C3177 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__conb_1_4/HI 0.00632f
C3178 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__inv_1_55/Y 2.51e-20
C3179 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_4/HI 0.00118f
C3180 sky130_fd_sc_hd__dfbbn_1_12/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00135f
C3181 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 8.55e-20
C3182 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 7.46e-20
C3183 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 6.4e-19
C3184 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 5.15e-19
C3185 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 4.94e-20
C3186 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 0.00596f
C3187 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# V_GND 6.62e-19
C3188 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 1.78e-19
C3189 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_581_47# 2.57e-19
C3190 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__conb_1_23/HI 2e-20
C3191 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0111f
C3192 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0011f
C3193 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# sky130_fd_sc_hd__inv_1_107/Y 2.99e-19
C3194 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/Q_N -9.56e-20
C3195 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# sky130_fd_sc_hd__nand3_1_2/Y 2.05e-21
C3196 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 0.0117f
C3197 sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__conb_1_31/HI 0.0377f
C3198 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.94e-19
C3199 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__conb_1_31/HI -0.00108f
C3200 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_1_57/Y 2.07e-19
C3201 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# V_GND -0.00299f
C3202 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 6.46e-19
C3203 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__conb_1_1/HI -3.03e-19
C3204 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 8.36e-20
C3205 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__conb_1_0/HI 9.48e-19
C3206 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# V_GND 1.81e-19
C3207 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# sky130_fd_sc_hd__inv_1_103/Y 3.75e-20
C3208 sky130_fd_sc_hd__dfbbn_1_30/Q_N FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00308f
C3209 sky130_fd_sc_hd__inv_1_19/Y sky130_fd_sc_hd__conb_1_12/HI 4.09e-22
C3210 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0228f
C3211 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# Reset 9.87e-19
C3212 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__conb_1_11/HI 0.00305f
C3213 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 0.0569f
C3214 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.014f
C3215 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__inv_1_56/Y 2.19e-20
C3216 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00144f
C3217 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__conb_1_42/HI 0.00451f
C3218 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 9.94e-19
C3219 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand2_8_3/Y 2.97e-19
C3220 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/Q_N -4.24e-20
C3221 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0409f
C3222 sky130_fd_sc_hd__inv_1_97/Y V_LOW 0.34f
C3223 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# Reset 3.96e-19
C3224 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 9.04e-19
C3225 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 1.2f
C3226 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.0378f
C3227 sky130_fd_sc_hd__inv_1_63/Y sky130_fd_sc_hd__conb_1_2/HI 5.75e-20
C3228 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__conb_1_2/HI 0.0012f
C3229 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.54e-21
C3230 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# -0.00375f
C3231 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__inv_1_102/Y 1.43e-19
C3232 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00494f
C3233 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.14e-20
C3234 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__conb_1_9/HI 1.02e-19
C3235 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 1.16e-19
C3236 FALLING_COUNTER.COUNT_SUB_DFF6.Q V_GND 0.965f
C3237 sky130_fd_sc_hd__nand2_1_4/a_113_47# V_GND -1.38e-20
C3238 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__inv_1_56/Y 5.54e-19
C3239 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 9.58e-21
C3240 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.24e-19
C3241 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 0.149f
C3242 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__conb_1_44/HI 0.149f
C3243 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__inv_1_55/Y 5.85e-22
C3244 sky130_fd_sc_hd__conb_1_1/LO Reset 0.00229f
C3245 sky130_fd_sc_hd__fill_4_87/VPB V_GND 0.424f
C3246 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# sky130_fd_sc_hd__inv_1_4/Y 7.05e-19
C3247 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 7.17e-21
C3248 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 1.76e-20
C3249 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 3.87e-20
C3250 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 1.4e-21
C3251 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__inv_1_20/Y 6.15e-19
C3252 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 3.39e-21
C3253 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 3.51e-21
C3254 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 1.86e-19
C3255 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00386f
C3256 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.92e-21
C3257 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_85/A 1.28e-20
C3258 sky130_fd_sc_hd__conb_1_26/HI V_GND 0.0709f
C3259 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 5.13e-19
C3260 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_16_0/Y 0.0108f
C3261 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 0.116f
C3262 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.14e-20
C3263 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00126f
C3264 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# sky130_fd_sc_hd__conb_1_5/HI 0.00484f
C3265 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.79e-19
C3266 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 1.31e-20
C3267 sky130_fd_sc_hd__dfbbn_1_18/Q_N FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0159f
C3268 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# 0.00203f
C3269 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.0102f
C3270 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.71e-21
C3271 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 9.96e-21
C3272 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 5.66e-20
C3273 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 2.16e-19
C3274 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 6.26e-21
C3275 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 9.83e-19
C3276 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 9.89e-20
C3277 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 0.00123f
C3278 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__conb_1_4/HI 8.88e-20
C3279 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__conb_1_42/HI -9.85e-19
C3280 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_1/LO 7.93e-20
C3281 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_2/A 0.0674f
C3282 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__inv_1_13/Y 2.08e-21
C3283 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 9.94e-20
C3284 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/Q_N 0.023f
C3285 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0302f
C3286 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_193_47# -0.0607f
C3287 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# 0.00117f
C3288 sky130_fd_sc_hd__inv_1_96/Y V_LOW 0.308f
C3289 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 0.192f
C3290 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__inv_1_18/Y 0.00764f
C3291 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# V_LOW 0.0205f
C3292 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__conb_1_23/HI 5.63e-21
C3293 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.45e-19
C3294 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_381_47# 2.64e-21
C3295 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 0.0012f
C3296 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 5.71e-20
C3297 sky130_fd_sc_hd__inv_1_10/Y sky130_fd_sc_hd__inv_16_2/Y 4.6e-21
C3298 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 5.71e-19
C3299 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_581_47# 5e-19
C3300 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# V_LOW -0.107f
C3301 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__inv_1_57/Y 2.22e-19
C3302 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# V_GND -0.0103f
C3303 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__conb_1_9/HI 0.00936f
C3304 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# -0.00381f
C3305 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__conb_1_36/HI -3.09e-19
C3306 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_6/HI 8.11e-21
C3307 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 2.45e-20
C3308 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# sky130_fd_sc_hd__conb_1_36/HI 4.35e-19
C3309 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_49/LO 6.63e-19
C3310 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 0.00242f
C3311 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 7.61e-20
C3312 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_8_3/Y 0.28f
C3313 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# 5.84e-19
C3314 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 2.92e-20
C3315 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# sky130_fd_sc_hd__inv_16_2/Y 0.0022f
C3316 sky130_fd_sc_hd__inv_1_99/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.107f
C3317 Reset FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00143f
C3318 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# sky130_fd_sc_hd__conb_1_11/HI -0.00236f
C3319 sky130_fd_sc_hd__inv_1_69/Y V_LOW 0.304f
C3320 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# V_LOW -0.0842f
C3321 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# V_GND 0.00756f
C3322 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_193_47# -0.0128f
C3323 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# V_LOW -0.321f
C3324 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# V_LOW 0.00672f
C3325 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__conb_1_45/HI -2.07e-19
C3326 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0714f
C3327 sky130_fd_sc_hd__inv_1_68/Y V_LOW 0.0288f
C3328 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# V_GND 0.00137f
C3329 sky130_fd_sc_hd__inv_1_20/Y V_GND -0.00328f
C3330 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_70/A 1.95e-19
C3331 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0423f
C3332 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__inv_1_10/Y 2.9e-19
C3333 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# V_GND -0.00502f
C3334 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__conb_1_13/HI 0.00188f
C3335 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# Reset 7.49e-21
C3336 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.41e-20
C3337 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 0.0416f
C3338 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_37/HI 3.92e-20
C3339 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 9.59e-21
C3340 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# -0.00141f
C3341 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.04e-19
C3342 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0.00392f
C3343 sky130_fd_sc_hd__inv_1_51/Y V_LOW 0.0305f
C3344 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0.0104f
C3345 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0.0112f
C3346 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 9.06e-20
C3347 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# V_GND 0.00412f
C3348 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# V_GND 0.0114f
C3349 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 4.89e-19
C3350 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# V_GND -0.00413f
C3351 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_16_2/Y 0.849f
C3352 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__inv_1_53/Y 0.00152f
C3353 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__inv_1_112/Y 4.94e-20
C3354 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# sky130_fd_sc_hd__inv_1_21/Y 0.00415f
C3355 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0532f
C3356 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_70/A 0.0591f
C3357 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00357f
C3358 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# 8.3e-21
C3359 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 6.82e-19
C3360 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# V_LOW -0.118f
C3361 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# V_GND 0.0211f
C3362 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_35/HI 1.62e-21
C3363 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__inv_1_107/Y 9.72e-20
C3364 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 2.6e-19
C3365 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.68e-19
C3366 sky130_fd_sc_hd__inv_1_70/A V_GND 0.129f
C3367 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# -2.53e-20
C3368 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 0.0354f
C3369 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 5.48e-19
C3370 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# Reset 0.0411f
C3371 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 1.71e-20
C3372 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_106/Y 5.11e-20
C3373 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_1_62/Y 5.21e-19
C3374 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__inv_1_101/Y 5.88e-19
C3375 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 3.49e-19
C3376 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 4.66e-19
C3377 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 0.00122f
C3378 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 5.05e-19
C3379 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0.00106f
C3380 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 9.94e-19
C3381 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# V_GND 0.0239f
C3382 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# V_GND 0.0127f
C3383 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0406f
C3384 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.91e-21
C3385 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 1.41e-20
C3386 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 1.5e-19
C3387 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# 1.72e-20
C3388 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__conb_1_4/HI 7.43e-21
C3389 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__conb_1_42/HI -2.07e-19
C3390 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_76/A 0.174f
C3391 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__conb_1_16/HI 0.105f
C3392 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# V_GND 0.00862f
C3393 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 1.29e-19
C3394 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_93/A 0.00619f
C3395 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# V_GND -0.00542f
C3396 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# 3.37e-19
C3397 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# V_LOW 9.28e-19
C3398 sky130_fd_sc_hd__nand2_1_0/a_113_47# V_LOW -1.78e-19
C3399 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# 2.43e-19
C3400 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 4.2e-19
C3401 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# sky130_fd_sc_hd__inv_1_60/Y 8.17e-19
C3402 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# V_LOW -0.00121f
C3403 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# -0.193f
C3404 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# V_LOW -2.09e-19
C3405 sky130_fd_sc_hd__dfbbn_1_20/Q_N RISING_COUNTER.COUNT_SUB_DFF1.Q 2.31e-19
C3406 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# -0.00141f
C3407 sky130_fd_sc_hd__inv_1_27/Y V_GND 0.118f
C3408 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__conb_1_36/HI -2.07e-19
C3409 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# V_LOW -0.103f
C3410 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# V_GND -0.145f
C3411 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# 7.35e-20
C3412 sky130_fd_sc_hd__inv_1_40/A V_LOW 0.0341f
C3413 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.33e-19
C3414 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 3.63e-19
C3415 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 8.95e-21
C3416 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# V_LOW -2.68e-19
C3417 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# V_GND -7.03e-19
C3418 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 0.00263f
C3419 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 2.67e-19
C3420 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# V_GND 9.12e-19
C3421 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.18e-20
C3422 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# -2.18e-19
C3423 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__nand3_1_1/Y 0.00209f
C3424 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# -5.54e-21
C3425 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.0133f
C3426 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# V_GND 0.00164f
C3427 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 3.56e-19
C3428 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 4.3e-21
C3429 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 6.46e-20
C3430 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00226f
C3431 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 8.74e-21
C3432 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_9/Y 1.57e-19
C3433 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# V_GND -4.22e-19
C3434 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# sky130_fd_sc_hd__conb_1_13/HI -0.00144f
C3435 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# V_LOW 3.56e-20
C3436 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__conb_1_41/HI 2.43e-20
C3437 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# -4.1e-19
C3438 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_891_329# -2.2e-20
C3439 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -6.43e-19
C3440 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# -0.0225f
C3441 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# sky130_fd_sc_hd__conb_1_37/HI 6.22e-22
C3442 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 2.76e-20
C3443 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_75/Y 0.00373f
C3444 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# V_GND 0.00159f
C3445 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.00292f
C3446 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# V_GND 0.00279f
C3447 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 5.28e-19
C3448 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 2.74e-19
C3449 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 4.97e-20
C3450 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 5.87e-20
C3451 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_891_329# 0.00134f
C3452 sky130_fd_sc_hd__inv_1_70/A sky130_fd_sc_hd__nand3_1_1/Y 7.96e-19
C3453 sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_1_63/Y 3.3e-19
C3454 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# V_GND 1.36e-19
C3455 sky130_fd_sc_hd__conb_1_16/LO V_GND -0.00524f
C3456 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# V_GND 2.4e-19
C3457 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# V_LOW 3.56e-20
C3458 sky130_fd_sc_hd__nand3_1_2/a_193_47# V_GND 8.56e-20
C3459 sky130_fd_sc_hd__conb_1_23/LO V_GND -0.00549f
C3460 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_473_413# 0.00646f
C3461 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_44/HI -0.00907f
C3462 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# V_LOW 2.26e-20
C3463 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 1.88e-19
C3464 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# V_GND -0.00521f
C3465 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# sky130_fd_sc_hd__inv_1_112/Y 8.08e-21
C3466 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# V_LOW -0.00121f
C3467 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/Q_N 9.27e-20
C3468 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.61e-20
C3469 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 7.48e-20
C3470 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# V_LOW -9.94e-19
C3471 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# V_GND 2.23e-19
C3472 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.98e-21
C3473 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# Reset 6.22e-19
C3474 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# V_GND -0.182f
C3475 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__conb_1_41/HI 1.02e-19
C3476 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# -1.44e-20
C3477 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_50/A 0.79f
C3478 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_381_47# -0.00175f
C3479 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__dfbbn_1_20/a_941_21# -6.22e-19
C3480 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# -0.00125f
C3481 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# Reset 2.59e-19
C3482 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 1.09e-20
C3483 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_95/A 3.98e-21
C3484 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 4.17e-20
C3485 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# V_GND 1.61e-19
C3486 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# 0.00715f
C3487 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.571f
C3488 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# V_GND 0.00189f
C3489 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00291f
C3490 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/Q_N 6.81e-21
C3491 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# -3.79e-20
C3492 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# -0.00336f
C3493 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# V_GND 0.00203f
C3494 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__inv_1_76/A 5.39e-21
C3495 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__conb_1_21/HI 0.00113f
C3496 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.024f
C3497 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# V_LOW -9.15e-19
C3498 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.59e-19
C3499 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# V_GND -3.75e-19
C3500 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__inv_1_54/Y 6.44e-19
C3501 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0.0149f
C3502 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 7.03e-19
C3503 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 3.52e-19
C3504 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 3.52e-19
C3505 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 7.03e-19
C3506 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 0.0149f
C3507 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00303f
C3508 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00642f
C3509 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.1e-20
C3510 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_46/HI 0.34f
C3511 sky130_fd_sc_hd__inv_1_107/Y sky130_fd_sc_hd__inv_16_1/Y 0.0345f
C3512 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_35/LO 0.0085f
C3513 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0458f
C3514 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_193_47# -0.0752f
C3515 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0288f
C3516 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.42e-19
C3517 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 1.93e-19
C3518 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 1.93e-19
C3519 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.0713f
C3520 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_26/HI 2.34e-19
C3521 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 5.18e-20
C3522 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__conb_1_44/HI 0.00752f
C3523 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# V_LOW -9.94e-19
C3524 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# V_LOW 4.8e-20
C3525 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# V_GND 1.08e-19
C3526 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.98e-19
C3527 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_15/Y 4.56e-21
C3528 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 1.49e-20
C3529 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# sky130_fd_sc_hd__inv_1_12/Y 2.45e-19
C3530 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__inv_1_65/Y 1.31e-20
C3531 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 3.38e-22
C3532 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 3.63e-20
C3533 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 3.68e-19
C3534 sky130_fd_sc_hd__conb_1_33/HI CLOCK_GEN.SR_Op.Q 2.8e-19
C3535 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__inv_1_12/Y 0.00104f
C3536 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.53e-20
C3537 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_1/Y 0.0227f
C3538 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.01e-19
C3539 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_63/Y 3.36e-20
C3540 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nand2_1_0/Y 0.0171f
C3541 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# V_LOW 0.0207f
C3542 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_381_47# 0.00171f
C3543 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_43/A 5.46e-20
C3544 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF3.Q 0.141f
C3545 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0025f
C3546 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_381_47# 0.0168f
C3547 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# V_LOW 0.00609f
C3548 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.75e-20
C3549 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__inv_1_10/Y 5.85e-22
C3550 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_41/HI -0.0135f
C3551 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# 2.84e-32
C3552 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# -0.00385f
C3553 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# -6.8e-19
C3554 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__conb_1_32/HI 0.00302f
C3555 sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# V_GND 1.4e-19
C3556 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# V_LOW -9.15e-19
C3557 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# V_GND -8.07e-19
C3558 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0137f
C3559 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# sky130_fd_sc_hd__conb_1_13/HI 5.19e-20
C3560 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 2.81e-20
C3561 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 7.26e-21
C3562 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00307f
C3563 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.93e-19
C3564 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 1.77e-20
C3565 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 7.13e-20
C3566 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 0.00144f
C3567 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# -5.33e-20
C3568 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_557_413# -3.67e-20
C3569 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.0457f
C3570 sky130_fd_sc_hd__inv_1_75/A sky130_fd_sc_hd__inv_1_80/A 2.37e-19
C3571 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.53e-21
C3572 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# 1.49e-19
C3573 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__conb_1_44/HI -9.71e-19
C3574 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.56e-20
C3575 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.1e-19
C3576 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# V_GND 0.00834f
C3577 sky130_fd_sc_hd__dfbbn_1_8/Q_N V_GND -0.0079f
C3578 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# V_GND 4.08e-19
C3579 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.5e-21
C3580 sky130_fd_sc_hd__conb_1_3/LO V_LOW 0.0728f
C3581 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 9.67e-19
C3582 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 5.52e-19
C3583 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.00391f
C3584 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 7.8e-19
C3585 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# V_GND 1.64e-19
C3586 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_94/A 0.295f
C3587 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_891_329# 0.00134f
C3588 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 5.36e-20
C3589 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# -2.37e-19
C3590 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_941_21# -0.00147f
C3591 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.00114f
C3592 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 4.03e-19
C3593 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0.0116f
C3594 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00278f
C3595 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.0116f
C3596 sky130_fd_sc_hd__conb_1_38/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.9e-20
C3597 sky130_fd_sc_hd__conb_1_27/LO V_LOW 0.0312f
C3598 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 4.14e-19
C3599 sky130_fd_sc_hd__conb_1_27/HI V_GND 0.269f
C3600 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__inv_1_98/Y 0.00104f
C3601 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# -6.29e-19
C3602 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_557_413# -3.67e-20
C3603 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# V_GND 0.00743f
C3604 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__conb_1_51/HI 0.0111f
C3605 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.021f
C3606 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 0.00256f
C3607 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# -4.66e-20
C3608 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# -3.79e-20
C3609 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_76/A 0.0161f
C3610 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.00121f
C3611 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 2.69e-21
C3612 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 1.75e-19
C3613 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 5.12e-20
C3614 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.29e-21
C3615 sky130_fd_sc_hd__inv_1_110/Y FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00171f
C3616 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__nand3_1_2/B 1.64e-20
C3617 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__inv_1_12/Y 0.0128f
C3618 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.0888f
C3619 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.00912f
C3620 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# -0.00336f
C3621 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# -3.79e-20
C3622 sky130_fd_sc_hd__conb_1_38/LO V_LOW 0.0927f
C3623 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 6.12e-19
C3624 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 6.12e-19
C3625 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 1.31e-19
C3626 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 9.54e-21
C3627 sky130_fd_sc_hd__inv_1_23/Y V_GND 0.0899f
C3628 sky130_fd_sc_hd__conb_1_43/HI FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0212f
C3629 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 8e-21
C3630 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 3.67e-21
C3631 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 3.83e-20
C3632 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# V_LOW 0.00141f
C3633 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 5.7e-19
C3634 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.298f
C3635 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 5.7e-19
C3636 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# -0.00115f
C3637 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 1.47e-20
C3638 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__conb_1_44/HI 1.22e-20
C3639 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0405f
C3640 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_11/LO 9.17e-19
C3641 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__conb_1_49/HI 4.28e-21
C3642 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.149f
C3643 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.0257f
C3644 RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.414f
C3645 Reset V_SENSE 0.168f
C3646 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.137f
C3647 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# V_LOW 0.0168f
C3648 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 3.25e-20
C3649 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# V_GND 0.0103f
C3650 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0333f
C3651 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_791_47# 8.28e-22
C3652 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 1.27e-21
C3653 sky130_fd_sc_hd__conb_1_8/HI V_LOW 0.125f
C3654 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 0.032f
C3655 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# V_LOW -6.55e-19
C3656 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# -2.65e-20
C3657 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/Q_N -4.24e-20
C3658 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 8.92e-19
C3659 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__inv_1_53/Y 0.00129f
C3660 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__conb_1_12/HI 0.034f
C3661 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# V_GND -0.00509f
C3662 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 3.45e-19
C3663 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_13/LO 7.5e-19
C3664 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__inv_1_21/Y 0.144f
C3665 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# sky130_fd_sc_hd__conb_1_32/HI 1.76e-19
C3666 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# V_GND 0.0039f
C3667 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# V_GND 0.00847f
C3668 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 0.00182f
C3669 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 0.00903f
C3670 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 5.56e-19
C3671 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0.00182f
C3672 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 5.56e-19
C3673 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0.00903f
C3674 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__inv_1_15/Y 0.00307f
C3675 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.34e-20
C3676 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 4.84e-19
C3677 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 4.13e-20
C3678 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF1.Q 3.25e-19
C3679 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_1_103/Y 0.00735f
C3680 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__conb_1_44/HI 4.59e-21
C3681 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# V_GND 8.28e-19
C3682 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_1_108/Y 0.00769f
C3683 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__conb_1_11/HI 2.57e-19
C3684 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__conb_1_27/HI 0.00591f
C3685 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_557_413# -0.0012f
C3686 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_891_329# -2.46e-19
C3687 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# -0.00946f
C3688 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# V_LOW 2.26e-20
C3689 sky130_fd_sc_hd__conb_1_44/LO V_GND -0.00517f
C3690 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 9.88e-20
C3691 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.3e-21
C3692 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0234f
C3693 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 5.43e-19
C3694 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_45/HI 0.0287f
C3695 CLOCK_GEN.SR_Op.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00267f
C3696 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 1.29e-21
C3697 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.5e-19
C3698 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF18.Q 0.105f
C3699 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__inv_16_1/Y 1.12e-19
C3700 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.87e-20
C3701 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# -7.17e-20
C3702 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# -1.66e-19
C3703 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/Q_N -9.56e-20
C3704 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0278f
C3705 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__conb_1_48/LO 1.88e-19
C3706 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 9.03e-19
C3707 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__inv_1_23/Y 2.39e-19
C3708 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0456f
C3709 sky130_fd_sc_hd__inv_1_11/Y V_GND 0.0967f
C3710 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__conb_1_8/HI 3.97e-20
C3711 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 5.04e-21
C3712 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00131f
C3713 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.87f
C3714 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# V_GND -0.00461f
C3715 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__conb_1_34/HI 4.02e-21
C3716 sky130_fd_sc_hd__dfbbn_1_50/a_1159_47# sky130_fd_sc_hd__conb_1_51/HI 8.86e-20
C3717 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# 7.25e-22
C3718 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0315f
C3719 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 8.22e-23
C3720 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 0.00128f
C3721 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 4.07e-21
C3722 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 2.16e-19
C3723 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 3.97e-20
C3724 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 8.77e-20
C3725 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 5.27e-20
C3726 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0.0113f
C3727 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.00174f
C3728 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# V_LOW 2.26e-20
C3729 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 0.00532f
C3730 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# sky130_fd_sc_hd__inv_1_12/Y 7.13e-19
C3731 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 0.0475f
C3732 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.3e-20
C3733 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.47e-20
C3734 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.404f
C3735 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_23/LO 0.00968f
C3736 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 0.00111f
C3737 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.169f
C3738 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 4.77e-20
C3739 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 1.92e-19
C3740 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/Q_N 1.98e-19
C3741 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_23/HI 2.54e-19
C3742 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 1.98e-19
C3743 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 6.61e-19
C3744 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.03f
C3745 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.00174f
C3746 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_71/Y 4.47e-20
C3747 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 5.7e-19
C3748 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.57e-21
C3749 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 2.59e-20
C3750 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.78e-20
C3751 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 4.72e-20
C3752 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 7.68e-19
C3753 FALLING_COUNTER.COUNT_SUB_DFF7.Q V_GND 0.759f
C3754 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.0018f
C3755 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 5.48e-21
C3756 sky130_fd_sc_hd__conb_1_22/HI V_GND 0.432f
C3757 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__conb_1_2/HI 0.0114f
C3758 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0271f
C3759 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00228f
C3760 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_581_47# -7.91e-19
C3761 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 8.44e-20
C3762 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_1_103/Y 0.0132f
C3763 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__conb_1_44/HI 4.28e-21
C3764 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# V_LOW 4.8e-20
C3765 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_106/Y 2.55e-21
C3766 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_16_1/Y 9.79e-19
C3767 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# V_GND 0.00319f
C3768 FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_15/Y 0.0176f
C3769 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 1.11f
C3770 sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__inv_1_97/Y 1.25e-19
C3771 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_119/Y 3.88e-19
C3772 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 6.55e-20
C3773 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 7.96e-19
C3774 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 3.26e-19
C3775 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# 5.02e-19
C3776 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_473_413# 0.0248f
C3777 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 7.56e-19
C3778 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.4e-20
C3779 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.00358f
C3780 sky130_fd_sc_hd__dfbbn_1_46/Q_N V_LOW -4.42e-19
C3781 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.54e-21
C3782 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 4.99e-19
C3783 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 2.83e-21
C3784 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 1.11e-20
C3785 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.62e-22
C3786 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# V_GND -0.00711f
C3787 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_78/A 0.0608f
C3788 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0.00103f
C3789 sky130_fd_sc_hd__conb_1_36/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.157f
C3790 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_17/Y 3.79e-19
C3791 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# V_GND 2.29e-19
C3792 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -1.89e-19
C3793 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# -2.52e-19
C3794 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.0427f
C3795 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.52e-21
C3796 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_54/Y 2.76e-21
C3797 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# V_GND 3.34e-19
C3798 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_647_21# 8.7e-21
C3799 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_791_47# 3.86e-19
C3800 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 3.86e-19
C3801 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0352f
C3802 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__inv_1_15/Y 1.46e-19
C3803 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_1_1/a_113_47# 1.89e-19
C3804 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_891_329# 6.98e-19
C3805 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 7.03e-19
C3806 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 7.03e-19
C3807 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# sky130_fd_sc_hd__inv_1_103/Y 2.67e-19
C3808 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 8.84e-20
C3809 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# sky130_fd_sc_hd__inv_1_108/Y 5.98e-19
C3810 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__conb_1_27/HI 0.00297f
C3811 sky130_fd_sc_hd__nand2_8_2/a_27_47# V_GND 2.8e-19
C3812 sky130_fd_sc_hd__fill_4_60/VPB V_LOW 0.797f
C3813 sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__inv_2_0/Y 4.5e-19
C3814 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# V_GND 0.00426f
C3815 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_891_329# -2.46e-19
C3816 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_557_413# -0.0012f
C3817 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# -0.00157f
C3818 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_1_47/Y 3.36e-20
C3819 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 1.34e-19
C3820 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__conb_1_35/HI 0.00211f
C3821 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 3.23e-20
C3822 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0205f
C3823 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# sky130_fd_sc_hd__inv_16_1/Y 2.27e-19
C3824 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0186f
C3825 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0302f
C3826 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 2.34e-20
C3827 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 3.52e-20
C3828 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.49e-20
C3829 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.24e-20
C3830 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_39/LO 0.00328f
C3831 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# sky130_fd_sc_hd__inv_1_23/Y 5.8e-19
C3832 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.73e-19
C3833 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.56e-21
C3834 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00113f
C3835 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__conb_1_0/HI 1.99e-19
C3836 sky130_fd_sc_hd__conb_1_17/LO V_LOW 0.0864f
C3837 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 3.35e-19
C3838 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.86e-20
C3839 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_27_47# 0.00125f
C3840 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 1.43e-21
C3841 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__inv_16_2/Y 8.98e-19
C3842 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.91e-20
C3843 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 3e-20
C3844 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 9.29e-21
C3845 sky130_fd_sc_hd__inv_1_107/Y V_LOW 0.0237f
C3846 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0223f
C3847 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.32e-21
C3848 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.089f
C3849 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_16_1/Y 0.00182f
C3850 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00655f
C3851 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 8.55e-20
C3852 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__conb_1_33/HI 6.53e-19
C3853 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 0.00317f
C3854 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00147f
C3855 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# -2.52e-19
C3856 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -3.88e-19
C3857 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# sky130_fd_sc_hd__inv_1_103/Y 2.47e-19
C3858 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 1.22e-21
C3859 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.0016f
C3860 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__inv_16_1/Y 0.0297f
C3861 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 9.79e-22
C3862 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 0.0255f
C3863 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# sky130_fd_sc_hd__conb_1_47/HI 1.44e-19
C3864 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 4.51e-19
C3865 sky130_fd_sc_hd__conb_1_50/HI V_GND 0.0527f
C3866 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_40/LO 1.47e-20
C3867 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# 7.6e-19
C3868 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 1.32e-20
C3869 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.33e-20
C3870 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# 5.07e-19
C3871 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# V_LOW 0.00606f
C3872 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 8.11e-21
C3873 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# V_LOW -0.104f
C3874 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.0101f
C3875 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 8.79e-22
C3876 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# V_LOW 4.8e-20
C3877 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00104f
C3878 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# V_LOW 0.0119f
C3879 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 1.32e-20
C3880 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# -4.98e-19
C3881 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# -0.0103f
C3882 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 8.71e-20
C3883 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_100/Y 0.0608f
C3884 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0555f
C3885 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.0397f
C3886 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# V_LOW 6.57e-19
C3887 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_16_1/Y 1.83e-20
C3888 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 2.38e-20
C3889 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 0.00123f
C3890 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_891_329# 3.21e-19
C3891 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# -1.76e-19
C3892 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 3.53e-19
C3893 sky130_fd_sc_hd__inv_1_28/Y V_SENSE 0.105f
C3894 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_91/A 0.0998f
C3895 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_119/Y -5.45e-20
C3896 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# V_LOW 0.00537f
C3897 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.0012f
C3898 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__inv_1_50/Y 5.11e-19
C3899 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# V_GND 3.37e-19
C3900 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# V_GND -0.00532f
C3901 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# V_LOW 0.00734f
C3902 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_381_47# 0.0145f
C3903 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# -6.23e-21
C3904 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_381_47# -4.5e-20
C3905 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 0.0305f
C3906 sky130_fd_sc_hd__dfbbn_1_15/a_581_47# V_GND 2.02e-19
C3907 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# V_GND 0.00157f
C3908 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# -4.36e-19
C3909 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# 1.23e-19
C3910 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# V_GND 2.6e-19
C3911 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# -0.00458f
C3912 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_647_21# -0.00431f
C3913 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 3.47e-21
C3914 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_2/HI 4.73e-19
C3915 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_647_21# -0.00431f
C3916 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_473_413# -0.00554f
C3917 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_941_21# 0.00343f
C3918 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_39/LO 0.00508f
C3919 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__conb_1_49/HI 0.0215f
C3920 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# sky130_fd_sc_hd__conb_1_0/HI 1.62e-19
C3921 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# V_GND 3.42e-19
C3922 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_15/LO 0.0124f
C3923 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0396f
C3924 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_1_59/Y 0.0106f
C3925 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# V_GND 0.0023f
C3926 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__conb_1_21/HI 4.13e-21
C3927 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# Reset 8.49e-19
C3928 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.13e-19
C3929 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0324f
C3930 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 8.52e-19
C3931 sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.52e-19
C3932 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# V_LOW 0.00126f
C3933 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# V_GND 0.0037f
C3934 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 1.91e-19
C3935 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.06e-19
C3936 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 1.68e-19
C3937 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_16_1/Y 5.11e-20
C3938 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.01e-20
C3939 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__inv_1_6/Y 6.34e-19
C3940 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.26e-20
C3941 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# -1.76e-19
C3942 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.116f
C3943 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_473_413# -0.00834f
C3944 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -1.61e-19
C3945 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 8.07e-20
C3946 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 1.15e-19
C3947 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 0.0119f
C3948 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00837f
C3949 FALLING_COUNTER.COUNT_SUB_DFF5.Q Reset 2.66f
C3950 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_95/A 0.115f
C3951 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_94/A 2.45e-19
C3952 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__inv_1_62/Y 0.00311f
C3953 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# -0.00813f
C3954 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__inv_16_0/Y 4.95e-19
C3955 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# V_GND 3.81e-19
C3956 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# sky130_fd_sc_hd__inv_1_11/Y 3.95e-19
C3957 sky130_fd_sc_hd__conb_1_20/HI V_LOW 0.13f
C3958 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# 3.29e-20
C3959 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 4.73e-21
C3960 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 6.84e-19
C3961 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# V_LOW -2.78e-35
C3962 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# V_LOW -9.94e-19
C3963 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 0.0118f
C3964 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_94/Y 0.0572f
C3965 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_8/HI 3.95e-20
C3966 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 2.44e-20
C3967 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 5.84e-21
C3968 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 2.26e-19
C3969 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_67/Y 1.42e-20
C3970 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 5.45e-20
C3971 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# V_LOW 1.79e-20
C3972 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 2.14e-19
C3973 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# -6.8e-19
C3974 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 4.04e-20
C3975 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 6.98e-19
C3976 sky130_fd_sc_hd__conb_1_10/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00122f
C3977 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 6.74e-19
C3978 sky130_fd_sc_hd__conb_1_26/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 9.84e-20
C3979 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# V_LOW -0.0502f
C3980 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_8_3/Y 0.0132f
C3981 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 1.94e-19
C3982 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_16_1/Y 0.157f
C3983 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__inv_1_102/Y 2.74e-19
C3984 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__conb_1_50/LO 1.33e-19
C3985 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_5/a_891_329# 3.48e-21
C3986 sky130_fd_sc_hd__conb_1_40/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 8.85e-20
C3987 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__nand2_8_0/a_27_47# 4.05e-20
C3988 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__inv_1_108/Y 1.17e-19
C3989 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__conb_1_13/HI 3.13e-20
C3990 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 0.0255f
C3991 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_22/HI 0.0419f
C3992 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0448f
C3993 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_15/HI 0.0014f
C3994 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.373f
C3995 FULL_COUNTER.COUNT_SUB_DFF4.Q V_GND 4.74f
C3996 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# V_LOW -2.78e-35
C3997 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0182f
C3998 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# V_GND -3.69e-19
C3999 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__conb_1_21/HI 0.0196f
C4000 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__inv_1_49/Y 0.035f
C4001 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_1_105/Y 9.13e-21
C4002 sky130_fd_sc_hd__nand2_8_5/a_27_47# V_GND -0.0569f
C4003 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0311f
C4004 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 3.37e-19
C4005 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# V_GND -0.169f
C4006 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 1.03e-20
C4007 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# V_GND 1.48e-19
C4008 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_21/HI 1.99e-19
C4009 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 4.74e-20
C4010 sky130_fd_sc_hd__conb_1_40/LO V_LOW 0.0955f
C4011 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# V_LOW 4.8e-20
C4012 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_93/A 2.21e-19
C4013 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 0.00103f
C4014 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# V_GND 0.00178f
C4015 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# CLOCK_GEN.SR_Op.Q 6.5e-19
C4016 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.0295f
C4017 FULL_COUNTER.COUNT_SUB_DFF7.Q V_GND 4.18f
C4018 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 9.87e-19
C4019 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.00139f
C4020 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.00108f
C4021 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__conb_1_46/HI 2.15e-20
C4022 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.0043f
C4023 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0012f
C4024 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.04e-19
C4025 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_193_47# -0.0508f
C4026 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# 7.25e-22
C4027 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.0137f
C4028 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 0.369f
C4029 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.59e-20
C4030 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# sky130_fd_sc_hd__conb_1_49/HI 0.0111f
C4031 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 9.42e-20
C4032 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# sky130_fd_sc_hd__inv_1_59/Y 7.18e-21
C4033 sky130_fd_sc_hd__conb_1_31/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0591f
C4034 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00475f
C4035 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# V_GND 0.00227f
C4036 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 1.58e-21
C4037 FULL_COUNTER.COUNT_SUB_DFF10.Q V_LOW 0.639f
C4038 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_891_329# 1.69e-21
C4039 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00267f
C4040 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.42e-19
C4041 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.68e-21
C4042 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00348f
C4043 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_891_329# 3.14e-19
C4044 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 1.72e-19
C4045 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# V_GND 0.0672f
C4046 sky130_fd_sc_hd__conb_1_51/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.3f
C4047 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0358f
C4048 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# -0.00813f
C4049 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# V_GND 2.05e-19
C4050 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# -3.79e-20
C4051 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# -4.66e-20
C4052 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 5.76e-20
C4053 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_20/HI 0.00741f
C4054 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 5.23e-22
C4055 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 5.23e-22
C4056 sky130_fd_sc_hd__inv_1_89/A Reset 0.0031f
C4057 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00405f
C4058 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 5.67e-19
C4059 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_86/Y 0.156f
C4060 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00358f
C4061 sky130_fd_sc_hd__conb_1_51/HI V_LOW 0.142f
C4062 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# -0.00149f
C4063 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0461f
C4064 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -0.0163f
C4065 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# -2.57e-20
C4066 FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_12/Y 1.17e-19
C4067 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/Q_N 9.37e-20
C4068 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 4.4e-19
C4069 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_647_21# 0.00692f
C4070 sky130_fd_sc_hd__inv_1_43/A V_GND 0.0526f
C4071 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# -5.54e-21
C4072 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_51/A 0.00228f
C4073 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_83/Y 0.0206f
C4074 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# -0.00141f
C4075 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00533f
C4076 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.0724f
C4077 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 4.61e-19
C4078 sky130_fd_sc_hd__conb_1_34/HI sky130_fd_sc_hd__inv_16_0/Y 0.0191f
C4079 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__inv_1_54/Y 2.04e-21
C4080 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# -0.00441f
C4081 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.05e-20
C4082 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 6.11e-19
C4083 sky130_fd_sc_hd__dfbbn_1_22/Q_N V_LOW 1.99e-19
C4084 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.24e-20
C4085 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_76/A 0.577f
C4086 sky130_fd_sc_hd__conb_1_41/HI sky130_fd_sc_hd__inv_16_1/Y 0.181f
C4087 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 0.0106f
C4088 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 7.21e-19
C4089 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_63/Y 0.0018f
C4090 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# V_LOW -9.15e-19
C4091 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 2.7e-21
C4092 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_381_47# -0.00869f
C4093 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 6.09e-19
C4094 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0294f
C4095 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00742f
C4096 sky130_fd_sc_hd__dfbbn_1_13/Q_N FULL_COUNTER.COUNT_SUB_DFF9.Q 1.83e-19
C4097 sky130_fd_sc_hd__dfbbn_1_39/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0323f
C4098 sky130_fd_sc_hd__dfbbn_1_45/Q_N V_LOW -0.00993f
C4099 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__inv_1_11/Y 0.00125f
C4100 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# V_LOW -2.68e-19
C4101 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.43e-20
C4102 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__inv_1_5/Y 1.31e-20
C4103 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__inv_16_0/Y 8.33e-21
C4104 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_50/A 0.0316f
C4105 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 9.66e-21
C4106 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 2.57e-22
C4107 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.27e-21
C4108 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.46e-21
C4109 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_15/HI 3.07e-19
C4110 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_1_90/Y 1.72e-20
C4111 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__conb_1_25/HI 0.00243f
C4112 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00826f
C4113 sky130_fd_sc_hd__dfbbn_1_18/Q_N V_LOW -7.65e-19
C4114 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__inv_1_9/Y 0.0131f
C4115 RISING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_60/Y 0.072f
C4116 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/Q_N -9.56e-20
C4117 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# V_GND 1.95e-19
C4118 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__conb_1_21/HI 1.62e-19
C4119 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 5.33e-21
C4120 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# V_LOW 1.85e-19
C4121 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# -4.66e-20
C4122 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# -3.79e-20
C4123 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 3.22e-21
C4124 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.4e-19
C4125 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__conb_1_37/HI -1.88e-20
C4126 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# CLOCK_GEN.SR_Op.Q 2.03e-19
C4127 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# 6.53e-19
C4128 sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# V_GND 1.36e-19
C4129 sky130_fd_sc_hd__dfbbn_1_24/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 0.00167f
C4130 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 3.9e-19
C4131 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 0.00114f
C4132 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__conb_1_30/HI 3.96e-19
C4133 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 8.11e-19
C4134 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 0.00188f
C4135 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 2.02e-20
C4136 FULL_COUNTER.COUNT_SUB_DFF19.Q V_LOW 1.57f
C4137 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.96e-19
C4138 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 3.16e-21
C4139 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 4.59e-21
C4140 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.72e-19
C4141 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 7.56e-21
C4142 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_45/A 1.59e-19
C4143 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 0.00188f
C4144 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__nand2_8_0/a_27_47# 4.25e-21
C4145 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 9.64e-20
C4146 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__conb_1_49/HI 0.00163f
C4147 sky130_fd_sc_hd__conb_1_38/HI FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00344f
C4148 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__inv_1_19/Y 0.00476f
C4149 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_891_329# 1.36e-19
C4150 sky130_fd_sc_hd__dfbbn_1_44/Q_N V_GND 0.0026f
C4151 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_44/A 0.038f
C4152 sky130_fd_sc_hd__conb_1_37/LO V_LOW 0.076f
C4153 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 8.48e-19
C4154 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 6.21e-21
C4155 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 7.37e-20
C4156 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 1.11e-20
C4157 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# V_GND 3.03e-19
C4158 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# -0.00107f
C4159 sky130_fd_sc_hd__dfbbn_1_25/Q_N V_LOW -0.0104f
C4160 sky130_fd_sc_hd__nand3_1_2/B sky130_fd_sc_hd__inv_1_67/Y 2.61e-20
C4161 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.01e-20
C4162 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_6/HI 0.00175f
C4163 sky130_fd_sc_hd__conb_1_48/LO V_LOW 0.0381f
C4164 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__conb_1_6/HI 0.0012f
C4165 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 6.35e-19
C4166 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 4.96e-19
C4167 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 3.39e-21
C4168 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__conb_1_37/LO 0.00469f
C4169 sky130_fd_sc_hd__conb_1_21/LO V_LOW 0.083f
C4170 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_581_47# -2.6e-20
C4171 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# -9.48e-19
C4172 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# CLOCK_GEN.SR_Op.Q 7.65e-21
C4173 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__inv_1_21/Y 0.253f
C4174 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_41/LO 1.19e-20
C4175 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 1.15e-19
C4176 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 1.97e-21
C4177 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.00523f
C4178 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 9.21e-20
C4179 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.01e-20
C4180 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00558f
C4181 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -3.34e-20
C4182 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 5.76e-20
C4183 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0058f
C4184 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 7.6e-20
C4185 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.19f
C4186 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# -0.00141f
C4187 sky130_fd_sc_hd__conb_1_15/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00127f
C4188 sky130_fd_sc_hd__dfbbn_1_13/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00399f
C4189 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# V_LOW -0.00298f
C4190 RISING_COUNTER.COUNT_SUB_DFF9.Q V_LOW 0.693f
C4191 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.104f
C4192 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.02e-20
C4193 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.34e-20
C4194 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# -0.00107f
C4195 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 7.27e-21
C4196 sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__inv_1_63/Y 1.69e-19
C4197 sky130_fd_sc_hd__inv_1_54/Y CLOCK_GEN.SR_Op.Q 0.423f
C4198 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.116f
C4199 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# 0.00193f
C4200 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# CLOCK_GEN.SR_Op.Q 5.04e-20
C4201 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00855f
C4202 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.22e-21
C4203 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 1.64f
C4204 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# CLOCK_GEN.SR_Op.Q 0.552f
C4205 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# V_LOW -0.317f
C4206 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_22/Y 0.0476f
C4207 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 1.15e-21
C4208 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 5.37e-20
C4209 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__nand3_1_0/Y 0.00168f
C4210 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 9.03e-19
C4211 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_76/A 2.63e-19
C4212 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 6.8e-21
C4213 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 5.59e-19
C4214 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0498f
C4215 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 2.95e-20
C4216 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# V_GND 3.32e-19
C4217 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00223f
C4218 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__conb_1_31/HI 2.42e-21
C4219 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 1.88e-20
C4220 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 1.17e-19
C4221 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__conb_1_26/HI 0.0156f
C4222 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_21/HI 0.13f
C4223 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/Q_N 5.03e-19
C4224 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 8.51e-20
C4225 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 1.8e-19
C4226 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0197f
C4227 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_119/Y 0.00707f
C4228 V_HIGH V_SENSE 0.724f
C4229 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 6.47e-22
C4230 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 8.58e-21
C4231 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_86/Y 0.108f
C4232 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__nand2_8_2/A 6.55e-20
C4233 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# V_GND 0.0202f
C4234 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 1.35e-19
C4235 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_6/Y 0.172f
C4236 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_112/Y 5.19e-20
C4237 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__inv_1_108/Y 3.01e-20
C4238 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__conb_1_42/HI 6.27e-19
C4239 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/Q_N 4.47e-19
C4240 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 0.0372f
C4241 sky130_fd_sc_hd__dfbbn_1_26/Q_N RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0292f
C4242 sky130_fd_sc_hd__inv_16_0/Y V_LOW 2.58f
C4243 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# sky130_fd_sc_hd__conb_1_6/HI 9.94e-22
C4244 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__nand3_1_2/B 0.241f
C4245 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__conb_1_21/HI 0.00884f
C4246 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 2.2e-20
C4247 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/Q_N 2.2e-20
C4248 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__conb_1_6/HI 5.99e-19
C4249 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 2.69e-21
C4250 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 9.29e-21
C4251 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 2.04e-21
C4252 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 5.99e-19
C4253 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.0033f
C4254 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 2.23e-20
C4255 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_85/Y 0.0212f
C4256 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_193_47# -0.0128f
C4257 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/Q_N 8.96e-21
C4258 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 9.91e-20
C4259 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__conb_1_16/HI 6.92e-20
C4260 Reset sky130_fd_sc_hd__inv_2_0/A 0.0245f
C4261 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/Q_N -4.33e-20
C4262 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_1_58/Y 1.85e-19
C4263 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI -0.0134f
C4264 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0556f
C4265 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.037f
C4266 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_16_1/Y 0.449f
C4267 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 4.56e-19
C4268 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 2.03e-20
C4269 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 4.02e-20
C4270 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# V_LOW -2.78e-35
C4271 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__conb_1_12/HI 2.41e-21
C4272 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_10/Q_N 1.31e-19
C4273 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 9.77e-21
C4274 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.95e-21
C4275 sky130_fd_sc_hd__inv_1_91/Y V_LOW 0.689f
C4276 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__conb_1_25/HI -0.00839f
C4277 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__conb_1_11/HI 1.5e-20
C4278 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00138f
C4279 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00576f
C4280 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__conb_1_2/HI 1.32e-20
C4281 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.0315f
C4282 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_26/Y 9.01e-20
C4283 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 6.77e-20
C4284 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# 0.0012f
C4285 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__conb_1_30/HI 0.00998f
C4286 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# -0.00108f
C4287 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.79e-19
C4288 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__conb_1_12/HI 6.82e-21
C4289 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# 4.67e-21
C4290 RISING_COUNTER.COUNT_SUB_DFF3.Q V_GND 1.49f
C4291 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.04e-20
C4292 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.03e-19
C4293 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_581_47# 3.74e-20
C4294 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00593f
C4295 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__inv_1_54/Y 0.00931f
C4296 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.88e-20
C4297 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_42/Y 0.0121f
C4298 sky130_fd_sc_hd__inv_1_39/Y V_LOW 0.141f
C4299 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_76/A 0.0382f
C4300 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 0.00696f
C4301 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 1.81e-19
C4302 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 6.33e-20
C4303 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00122f
C4304 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/Q_N -1.42e-32
C4305 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# V_LOW 0.0159f
C4306 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__conb_1_28/HI 9.87e-21
C4307 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# sky130_fd_sc_hd__conb_1_31/HI 1.5e-20
C4308 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.011f
C4309 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_94/Y 0.0214f
C4310 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_941_21# 0.0496f
C4311 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00408f
C4312 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__inv_16_0/Y -2.12e-19
C4313 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 1.02e-19
C4314 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# 1.92e-22
C4315 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0352f
C4316 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# -0.234f
C4317 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# V_GND 1.82e-19
C4318 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__conb_1_6/HI 5.57e-21
C4319 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 1.68e-19
C4320 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.607f
C4321 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00292f
C4322 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_473_413# -8.15e-19
C4323 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 0.00172f
C4324 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# CLOCK_GEN.SR_Op.Q 1.98e-20
C4325 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_22/HI 4.95e-20
C4326 sky130_fd_sc_hd__conb_1_43/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.15e-19
C4327 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# V_LOW 0.0135f
C4328 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_97/A 7.68e-19
C4329 sky130_fd_sc_hd__fill_4_58/VPB V_GND 0.396f
C4330 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# 4.53e-19
C4331 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_25/HI 1.16e-19
C4332 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 1.49e-19
C4333 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_49/HI 4.84e-20
C4334 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# V_GND -0.00565f
C4335 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0122f
C4336 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0196f
C4337 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# V_LOW 0.00484f
C4338 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 4.03e-21
C4339 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# V_LOW 0.0136f
C4340 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# V_GND -0.151f
C4341 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.86e-19
C4342 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__conb_1_21/HI 2.04e-19
C4343 FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_41/HI 5.23e-21
C4344 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_53/Y 4.48e-20
C4345 sky130_fd_sc_hd__inv_1_93/Y V_LOW 0.0345f
C4346 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 5.02e-19
C4347 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# -0.00375f
C4348 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_6/Y 0.00318f
C4349 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 1.65e-19
C4350 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.16e-19
C4351 sky130_fd_sc_hd__inv_1_4/Y V_GND 0.0483f
C4352 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_18/HI 0.0051f
C4353 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_5/HI 7.36e-19
C4354 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# sky130_fd_sc_hd__inv_1_98/Y 6.07e-20
C4355 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# V_GND 5.95e-19
C4356 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_18/HI 0.154f
C4357 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__conb_1_18/HI 0.0115f
C4358 sky130_fd_sc_hd__conb_1_41/HI V_LOW 0.181f
C4359 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# V_GND 0.00429f
C4360 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__conb_1_17/HI 1.22e-21
C4361 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00804f
C4362 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__conb_1_23/HI 0.00357f
C4363 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 1.32e-19
C4364 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0.0359f
C4365 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# V_GND 0.00504f
C4366 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.61e-20
C4367 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 3.01e-19
C4368 sky130_fd_sc_hd__dfbbn_1_39/Q_N V_LOW -0.00141f
C4369 RISING_COUNTER.COUNT_SUB_DFF13.Q V_GND 1.58f
C4370 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/Q_N 3.71e-20
C4371 sky130_fd_sc_hd__inv_1_81/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00151f
C4372 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__conb_1_28/HI 0.014f
C4373 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# 1.41e-19
C4374 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.06e-21
C4375 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# sky130_fd_sc_hd__conb_1_25/HI -9.41e-19
C4376 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__inv_1_106/Y 0.00115f
C4377 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_941_21# -5.77e-20
C4378 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# -2.52e-19
C4379 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# -0.0187f
C4380 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# 0.00107f
C4381 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 7.56e-19
C4382 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 5.86e-22
C4383 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_581_47# -2.6e-20
C4384 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_193_47# -0.156f
C4385 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__conb_1_51/HI 5.69e-20
C4386 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_10/HI 2.62e-19
C4387 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 0.0409f
C4388 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 1.55e-20
C4389 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 5.91e-21
C4390 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# V_GND -0.151f
C4391 RISING_COUNTER.COUNT_SUB_DFF1.Q CLOCK_GEN.SR_Op.Q 0.109f
C4392 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 4.12e-19
C4393 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.38e-19
C4394 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__conb_1_22/HI 0.0225f
C4395 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# V_GND -0.174f
C4396 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__conb_1_17/HI 0.0683f
C4397 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__inv_1_16/Y 0.0275f
C4398 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -0.00164f
C4399 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# -2.25e-19
C4400 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 2.84e-32
C4401 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 4.88e-19
C4402 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__conb_1_20/LO 0.0519f
C4403 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__conb_1_16/HI 0.00296f
C4404 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_1_18/Y 5.63e-20
C4405 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.12e-19
C4406 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# V_LOW 0.00734f
C4407 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# 6.67e-22
C4408 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_12/HI 2.33e-19
C4409 sky130_fd_sc_hd__inv_1_91/A V_GND 0.0863f
C4410 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.00265f
C4411 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# 0.00165f
C4412 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# V_LOW -9.15e-19
C4413 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/Q_N 2.24e-20
C4414 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 3.15e-20
C4415 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 4.03e-21
C4416 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.84e-20
C4417 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# sky130_fd_sc_hd__conb_1_6/HI -2.65e-20
C4418 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# V_GND 5.27e-19
C4419 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__inv_1_61/Y 0.003f
C4420 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00418f
C4421 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.17e-19
C4422 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_70/Y 0.00155f
C4423 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_39/HI -1.06e-19
C4424 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.03e-19
C4425 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 3.67e-21
C4426 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 8e-21
C4427 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_46/HI 2.35e-20
C4428 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# CLOCK_GEN.SR_Op.Q 4.96e-19
C4429 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# 2.09e-19
C4430 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.13e-20
C4431 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__inv_1_18/Y 0.0319f
C4432 sky130_fd_sc_hd__inv_1_86/Y V_LOW 0.0218f
C4433 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__conb_1_12/LO 1.56e-20
C4434 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# -1.62e-20
C4435 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# -3.69e-19
C4436 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 0.0167f
C4437 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.7e-19
C4438 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# sky130_fd_sc_hd__inv_1_57/Y 3.18e-19
C4439 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# V_GND 3.44e-19
C4440 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# V_GND 3.61e-19
C4441 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 2.26e-21
C4442 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__inv_1_99/Y 1.31e-20
C4443 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.021f
C4444 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# V_LOW 2.94e-20
C4445 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.83e-19
C4446 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_107/Y 0.0264f
C4447 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# V_LOW 2.94e-20
C4448 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__conb_1_35/HI 0.00137f
C4449 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# V_GND 9.69e-20
C4450 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 4.5e-19
C4451 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 9.57e-19
C4452 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# sky130_fd_sc_hd__conb_1_40/HI 5.03e-19
C4453 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 6.21e-20
C4454 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 9.44e-19
C4455 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 8.86e-20
C4456 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0325f
C4457 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# -0.00141f
C4458 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 1.65e-20
C4459 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 1.77e-20
C4460 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_9/HI 0.0294f
C4461 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__inv_1_6/Y 1.07e-21
C4462 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.6e-20
C4463 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__conb_1_44/HI 7.1e-19
C4464 sky130_fd_sc_hd__conb_1_17/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00258f
C4465 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.52e-20
C4466 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_68/A 2.27e-19
C4467 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# V_GND -0.0112f
C4468 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 4.74e-19
C4469 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__conb_1_18/HI 0.0174f
C4470 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__nand3_1_0/Y 7.27e-19
C4471 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# V_GND 6.75e-19
C4472 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__conb_1_38/HI -0.00274f
C4473 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# V_LOW 3.56e-20
C4474 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_1/HI 5.02e-21
C4475 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_27/Q_N 0.0216f
C4476 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# 6.41e-19
C4477 sky130_fd_sc_hd__dfbbn_1_50/a_1159_47# V_GND 0.0011f
C4478 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# V_LOW -9.15e-19
C4479 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 4.64e-19
C4480 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00442f
C4481 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_647_21# 5.83e-19
C4482 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# -2.65e-20
C4483 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_21/Y 2.41e-19
C4484 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__conb_1_45/HI 0.001f
C4485 sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__conb_1_12/HI 3.41e-19
C4486 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__dfbbn_1_47/Q_N -1.83e-19
C4487 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00294f
C4488 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_9/LO 1.39e-20
C4489 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__nor2_1_0/Y 4.96e-20
C4490 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0443f
C4491 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# -1.76e-19
C4492 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.22e-20
C4493 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_78/A 7.08e-21
C4494 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.87e-21
C4495 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_17/HI 0.344f
C4496 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# V_LOW -0.00266f
C4497 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# V_GND 1.53e-19
C4498 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 3.42e-20
C4499 sky130_fd_sc_hd__conb_1_2/LO V_GND 0.00426f
C4500 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# sky130_fd_sc_hd__conb_1_22/HI 4.96e-20
C4501 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# V_GND 1.23e-19
C4502 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# -7.17e-20
C4503 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.28e-20
C4504 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# -1.63e-19
C4505 sky130_fd_sc_hd__inv_16_1/Y V_GND 6.09f
C4506 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# sky130_fd_sc_hd__conb_1_16/HI 0.00161f
C4507 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 1.63e-20
C4508 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 8.84e-20
C4509 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 9.87e-21
C4510 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__conb_1_12/HI -2.07e-19
C4511 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# -3.65e-19
C4512 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# -3.07e-19
C4513 sky130_fd_sc_hd__dfbbn_1_48/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0406f
C4514 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 4.72e-19
C4515 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_40/HI 0.00393f
C4516 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_14/Y 6.95e-21
C4517 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_98/Y 0.00791f
C4518 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_106/Y 0.613f
C4519 sky130_fd_sc_hd__inv_1_110/Y FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.38f
C4520 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 2.66e-22
C4521 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_22/Y 2.25e-20
C4522 Reset sky130_fd_sc_hd__inv_1_5/Y 6.26e-19
C4523 sky130_fd_sc_hd__conb_1_24/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00953f
C4524 sky130_fd_sc_hd__conb_1_29/LO V_GND -0.00282f
C4525 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# V_GND -8.16e-19
C4526 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0593f
C4527 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00366f
C4528 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__conb_1_39/HI -0.00653f
C4529 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 3.7e-21
C4530 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00104f
C4531 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# -1.76e-19
C4532 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# 0.00142f
C4533 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# V_GND 0.00972f
C4534 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# V_GND 0.00501f
C4535 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0985f
C4536 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_891_329# -3.3e-20
C4537 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# -0.00913f
C4538 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00136f
C4539 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__conb_1_32/HI -4.51e-19
C4540 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.06e-19
C4541 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.57e-19
C4542 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# sky130_fd_sc_hd__conb_1_35/HI 0.00258f
C4543 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_83/Y 2.01e-19
C4544 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF10.Q 4.44e-19
C4545 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# -0.00543f
C4546 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# Reset 4.26e-20
C4547 sky130_fd_sc_hd__conb_1_19/HI V_GND 0.0279f
C4548 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 9.81e-21
C4549 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_27/LO 1.85e-21
C4550 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.85e-19
C4551 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_93/A 0.00597f
C4552 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_76/A 0.00212f
C4553 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__inv_1_103/Y 2.73e-19
C4554 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# -0.00149f
C4555 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_1_58/Y 0.00693f
C4556 sky130_fd_sc_hd__conb_1_39/HI V_LOW 0.04f
C4557 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.016f
C4558 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_35/HI 4.89e-19
C4559 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 4.4e-21
C4560 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__conb_1_18/HI 0.0292f
C4561 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_67/Y 2.11e-19
C4562 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# sky130_fd_sc_hd__conb_1_38/HI -8.94e-19
C4563 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# V_GND -0.00164f
C4564 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_11/LO 5.04e-21
C4565 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_12/LO 2.18e-19
C4566 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 1.23e-19
C4567 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_15/HI 1.82e-21
C4568 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__conb_1_42/HI 4.37e-19
C4569 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__inv_1_7/Y 1.72e-19
C4570 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_16_2/Y 0.106f
C4571 sky130_fd_sc_hd__inv_1_83/Y V_GND 0.842f
C4572 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_75/A 1.01f
C4573 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__conb_1_34/HI 8.8e-20
C4574 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_63/Y 0.00229f
C4575 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 8.23e-19
C4576 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 3.52e-20
C4577 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 6.43e-20
C4578 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# -0.00198f
C4579 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_891_329# -2.2e-20
C4580 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.13e-20
C4581 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/Q_N 0.019f
C4582 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.2e-21
C4583 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__conb_1_51/LO 1.31e-20
C4584 sky130_fd_sc_hd__conb_1_28/HI V_LOW 0.0321f
C4585 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 0.005f
C4586 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__conb_1_48/HI 1.28e-19
C4587 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__inv_1_55/Y 0.00882f
C4588 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__conb_1_16/HI -7.91e-20
C4589 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# -0.0195f
C4590 sky130_fd_sc_hd__inv_1_32/A V_GND 0.106f
C4591 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.21e-20
C4592 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# V_LOW -9.15e-19
C4593 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 4.09e-20
C4594 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# V_LOW 4.8e-20
C4595 sky130_fd_sc_hd__dfbbn_1_42/Q_N V_LOW -0.00121f
C4596 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0.00421f
C4597 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 3.77e-19
C4598 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 3.29e-19
C4599 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__inv_1_59/Y 0.00249f
C4600 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# -1.65e-19
C4601 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# -7.17e-20
C4602 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# 3.02e-19
C4603 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__inv_1_57/Y 0.0153f
C4604 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__conb_1_40/HI 5.84e-19
C4605 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0565f
C4606 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 4.41e-20
C4607 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 5.03e-19
C4608 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 5.03e-19
C4609 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 4.41e-20
C4610 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0828f
C4611 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.24e-19
C4612 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00219f
C4613 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_112/Y 1.15e-19
C4614 sky130_fd_sc_hd__conb_1_34/HI V_GND 0.0532f
C4615 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00885f
C4616 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0342f
C4617 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__inv_1_100/Y 2.34e-20
C4618 sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__conb_1_12/LO 9.43e-20
C4619 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 3.81e-19
C4620 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# V_GND 0.0322f
C4621 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 8.82e-20
C4622 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_381_47# 0.0141f
C4623 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0295f
C4624 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 8.92e-21
C4625 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# V_GND 1.95e-19
C4626 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# V_GND 2.44e-19
C4627 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.414f
C4628 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# 1.42e-32
C4629 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# -0.00592f
C4630 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# V_LOW 4.8e-20
C4631 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__conb_1_32/HI -8.72e-19
C4632 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_473_413# 0.00215f
C4633 sky130_fd_sc_hd__dfbbn_1_6/Q_N V_LOW -0.00461f
C4634 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# -0.00141f
C4635 sky130_fd_sc_hd__conb_1_31/LO V_GND -0.00636f
C4636 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__nand3_1_2/Y 3.99e-20
C4637 sky130_fd_sc_hd__nand3_1_1/a_193_47# sky130_fd_sc_hd__inv_1_71/Y 3.1e-19
C4638 sky130_fd_sc_hd__dfbbn_1_22/Q_N RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00373f
C4639 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__conb_1_0/HI 0.0117f
C4640 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# V_GND 3.26e-19
C4641 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__inv_1_103/Y 1.42e-19
C4642 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_581_47# -2.6e-20
C4643 sky130_fd_sc_hd__inv_1_64/Y Reset 0.00296f
C4644 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.00269f
C4645 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# Reset 0.0334f
C4646 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_18/LO 8.81e-20
C4647 sky130_fd_sc_hd__conb_1_42/LO V_GND -0.00456f
C4648 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_381_47# 4.36e-19
C4649 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_61/Y 0.0697f
C4650 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_13/Q_N 0.00125f
C4651 sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__conb_1_38/HI 6.47e-19
C4652 sky130_fd_sc_hd__dfbbn_1_24/a_581_47# V_GND 2.65e-19
C4653 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__conb_1_34/HI 0.00498f
C4654 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 1.58e-21
C4655 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_50/Y 0.0997f
C4656 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_16/HI 0.0383f
C4657 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_14/LO 0.0308f
C4658 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.78e-19
C4659 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00337f
C4660 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.552f
C4661 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.72e-20
C4662 sky130_fd_sc_hd__inv_1_72/Y Reset 1.55e-19
C4663 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_1_0/Y 0.0145f
C4664 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_891_329# -2.46e-19
C4665 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_557_413# -0.0012f
C4666 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# -0.00436f
C4667 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# 7.02e-21
C4668 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 7.26e-19
C4669 sky130_fd_sc_hd__dfbbn_1_45/Q_N FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.1e-21
C4670 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 5e-21
C4671 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# -0.00385f
C4672 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 1.3e-19
C4673 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__conb_1_9/HI 1.83e-19
C4674 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00611f
C4675 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 8.32e-19
C4676 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0.00127f
C4677 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# 5.06e-19
C4678 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# sky130_fd_sc_hd__conb_1_48/HI 3.64e-19
C4679 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__conb_1_5/LO 1.16e-20
C4680 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 1.5e-19
C4681 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# V_LOW -9.15e-19
C4682 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.012f
C4683 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_65/Y 1.16e-19
C4684 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0967f
C4685 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_43/A 0.0652f
C4686 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 0.00104f
C4687 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# sky130_fd_sc_hd__inv_1_57/Y 1.98e-19
C4688 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__inv_1_22/Y 2.58e-19
C4689 sky130_fd_sc_hd__conb_1_9/LO sky130_fd_sc_hd__inv_16_2/Y 0.00698f
C4690 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0141f
C4691 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 3.94e-19
C4692 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 3.94e-19
C4693 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.54e-20
C4694 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_1_60/Y 1.74e-19
C4695 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 1.54e-20
C4696 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__conb_1_5/HI 0.0171f
C4697 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_16_0/Y 0.00238f
C4698 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.33e-19
C4699 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.64e-19
C4700 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_31/A 0.194f
C4701 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 1.44e-19
C4702 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 9.22e-20
C4703 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 9.22e-20
C4704 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_65/Y 0.00417f
C4705 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0.0811f
C4706 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# V_LOW 7.71e-19
C4707 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# V_LOW 2.26e-20
C4708 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_381_47# 0.0128f
C4709 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00491f
C4710 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__conb_1_4/HI 3.7e-19
C4711 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 6.36e-21
C4712 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 7.23e-19
C4713 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# V_GND 1.05e-19
C4714 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 3.88e-19
C4715 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 9.08e-19
C4716 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 3.22e-19
C4717 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 0.00334f
C4718 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0.00401f
C4719 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_34/a_381_47# 2.9e-19
C4720 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 1.97e-20
C4721 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_71/Y 0.0119f
C4722 sky130_fd_sc_hd__conb_1_46/LO sky130_fd_sc_hd__inv_16_1/Y 0.0305f
C4723 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__conb_1_32/HI -1.82e-19
C4724 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# 0.002f
C4725 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_47/HI 0.0097f
C4726 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI 8.11e-21
C4727 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 1.37f
C4728 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# sky130_fd_sc_hd__inv_1_107/Y 8.05e-20
C4729 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__nand3_1_2/Y 6.08e-21
C4730 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0736f
C4731 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.9e-21
C4732 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 0.0254f
C4733 sky130_fd_sc_hd__conb_1_48/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.011f
C4734 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 2.37e-19
C4735 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# V_GND -0.00461f
C4736 sky130_fd_sc_hd__inv_1_64/A V_LOW 0.297f
C4737 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# sky130_fd_sc_hd__conb_1_0/HI 2.04e-19
C4738 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__conb_1_1/HI -0.00174f
C4739 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# V_GND -0.00489f
C4740 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 4.23e-20
C4741 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# sky130_fd_sc_hd__inv_1_103/Y 6.13e-21
C4742 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_16_1/Y 7.69e-19
C4743 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# sky130_fd_sc_hd__conb_1_36/HI 2.05e-19
C4744 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# Reset 0.00149f
C4745 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 4.06e-21
C4746 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_51/HI 0.0018f
C4747 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# sky130_fd_sc_hd__inv_1_61/Y 1.6e-20
C4748 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_11/HI 0.0215f
C4749 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# sky130_fd_sc_hd__conb_1_34/HI 2.09e-19
C4750 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00924f
C4751 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_42/HI 3.7e-19
C4752 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 0.00861f
C4753 FALLING_COUNTER.COUNT_SUB_DFF0.Q V_GND 1.72f
C4754 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_75/A 9.81e-20
C4755 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/Q_N -9.56e-20
C4756 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00245f
C4757 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__conb_1_38/HI 9.12e-19
C4758 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# Reset 4.11e-19
C4759 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00138f
C4760 sky130_fd_sc_hd__inv_1_66/Y V_LOW 0.144f
C4761 sky130_fd_sc_hd__conb_1_21/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 5.69e-19
C4762 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# -5.42e-19
C4763 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 0.0204f
C4764 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# sky130_fd_sc_hd__conb_1_2/HI 2.11e-19
C4765 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.78e-21
C4766 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_557_413# -0.0012f
C4767 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# -0.0306f
C4768 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__inv_1_102/Y 0.00921f
C4769 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0123f
C4770 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.8e-20
C4771 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_1_56/Y -5.28e-20
C4772 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_11/HI 0.00204f
C4773 V_GND V_LOW 0.224p
C4774 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 0.0178f
C4775 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 2.35e-21
C4776 sky130_fd_sc_hd__conb_1_13/HI V_GND -0.115f
C4777 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_21/Y 0.282f
C4778 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__inv_1_4/Y 3.75e-21
C4779 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 1.37e-20
C4780 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 6.87e-22
C4781 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 4.46e-20
C4782 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 2.97e-19
C4783 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 2.07e-19
C4784 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 1.44e-19
C4785 sky130_fd_sc_hd__inv_1_106/Y V_LOW 0.177f
C4786 sky130_fd_sc_hd__dfbbn_1_48/a_581_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00108f
C4787 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_76/A 0.0177f
C4788 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00127f
C4789 sky130_fd_sc_hd__conb_1_36/LO V_GND -0.00332f
C4790 sky130_fd_sc_hd__inv_1_59/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.237f
C4791 sky130_fd_sc_hd__inv_2_0/A V_HIGH 0.0641f
C4792 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_16_0/Y 0.327f
C4793 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.06e-20
C4794 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__inv_1_60/Y 2.18e-20
C4795 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 0.0333f
C4796 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.42e-20
C4797 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0177f
C4798 sky130_fd_sc_hd__dfbbn_1_19/a_581_47# sky130_fd_sc_hd__conb_1_5/HI 3.08e-19
C4799 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.58e-19
C4800 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 0.0419f
C4801 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 1.66e-19
C4802 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 1.66e-19
C4803 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# 4.48e-21
C4804 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 2.58e-20
C4805 sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__conb_1_30/HI 4.26e-19
C4806 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 9.68e-21
C4807 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 7.59e-20
C4808 sky130_fd_sc_hd__dfbbn_1_29/Q_N RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0253f
C4809 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 1.1e-20
C4810 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 3.23e-19
C4811 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 8.9e-21
C4812 sky130_fd_sc_hd__conb_1_47/LO V_GND 0.00327f
C4813 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__conb_1_42/HI -0.00852f
C4814 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# sky130_fd_sc_hd__conb_1_4/HI -2.65e-20
C4815 sky130_fd_sc_hd__inv_1_12/Y V_LOW 0.417f
C4816 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_10/LO 8.84e-20
C4817 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 5.85e-19
C4818 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__conb_1_44/HI 0.135f
C4819 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.286f
C4820 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_647_21# -1.69e-19
C4821 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# 6.89e-20
C4822 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_76/A 0.0405f
C4823 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_2_0/Y 4.79e-21
C4824 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_22/Y 0.103f
C4825 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q -2.71e-20
C4826 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0277f
C4827 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# V_LOW 0.00578f
C4828 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_32/HI 0.0503f
C4829 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 0.00555f
C4830 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1_76/A 7.7e-19
C4831 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.29e-19
C4832 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 9.31e-19
C4833 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 1.3e-19
C4834 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# 2.81e-19
C4835 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# V_LOW 0.00888f
C4836 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 6.07e-20
C4837 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__conb_1_31/HI 3.75e-20
C4838 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# V_GND -0.00534f
C4839 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# sky130_fd_sc_hd__conb_1_9/HI -0.0018f
C4840 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# sky130_fd_sc_hd__conb_1_10/HI 1.08e-19
C4841 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_557_413# -3.67e-20
C4842 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# -0.0238f
C4843 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# sky130_fd_sc_hd__conb_1_36/HI -0.00581f
C4844 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__conb_1_1/HI -2.07e-19
C4845 sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__inv_1_71/A 3.15e-19
C4846 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 0.081f
C4847 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_1_22/Y 1.59e-19
C4848 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 1.73e-19
C4849 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 2.13e-20
C4850 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# 1.46e-19
C4851 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 0.00295f
C4852 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__conb_1_51/HI 1e-19
C4853 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_3/HI 0.142f
C4854 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# V_LOW 0.00304f
C4855 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# V_GND 0.00767f
C4856 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# V_LOW -0.00229f
C4857 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# V_GND 0.0214f
C4858 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# -0.00108f
C4859 sky130_fd_sc_hd__nand3_1_1/Y V_LOW 0.256f
C4860 sky130_fd_sc_hd__dfbbn_1_7/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0058f
C4861 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# V_LOW 0.0157f
C4862 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__conb_1_6/HI 0.0362f
C4863 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 7.34e-20
C4864 sky130_fd_sc_hd__conb_1_22/LO sky130_fd_sc_hd__conb_1_22/HI 0.00338f
C4865 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# sky130_fd_sc_hd__conb_1_45/HI 0.00109f
C4866 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# V_GND 0.00385f
C4867 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.202f
C4868 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_58/Y 1.03e-20
C4869 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0172f
C4870 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__inv_1_10/Y 0.0107f
C4871 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# V_GND 2.09e-19
C4872 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__conb_1_9/LO 8.84e-20
C4873 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_13/HI 0.0149f
C4874 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# Reset 0.00159f
C4875 sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__inv_1_85/A 7.53e-21
C4876 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__inv_16_1/Y 0.00113f
C4877 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.65e-19
C4878 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 6.71e-20
C4879 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_15/HI 0.00721f
C4880 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_24/HI 1.31e-20
C4881 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_58/Y 5.28e-20
C4882 Reset sky130_fd_sc_hd__nand2_8_9/Y 0.0922f
C4883 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 9.85e-20
C4884 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 5.76e-19
C4885 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 9.66e-19
C4886 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__inv_1_108/Y 0.00126f
C4887 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# V_GND 3.06e-19
C4888 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# V_GND 0.00287f
C4889 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# V_GND -0.00485f
C4890 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00107f
C4891 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__inv_1_112/Y 0.0686f
C4892 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# sky130_fd_sc_hd__inv_1_21/Y 1.1e-19
C4893 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00114f
C4894 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_12/HI 6.8e-20
C4895 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0346f
C4896 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 7.8e-21
C4897 sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__inv_16_0/Y 0.624f
C4898 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 3.69e-19
C4899 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# V_LOW -0.0155f
C4900 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0462f
C4901 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# V_GND 0.00682f
C4902 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00218f
C4903 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__inv_1_107/Y 5.47e-19
C4904 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 6.49e-20
C4905 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_76/A 1.12e-19
C4906 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.55e-19
C4907 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0405f
C4908 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# -5.33e-20
C4909 sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__inv_1_86/Y 1.23e-20
C4910 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_557_413# -3.67e-20
C4911 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 7.69e-20
C4912 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0911f
C4913 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# Reset 0.0434f
C4914 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 1.18e-20
C4915 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_106/Y 2.33e-20
C4916 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_89/Y 0.121f
C4917 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__inv_1_62/Y 9.61e-20
C4918 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 0.0035f
C4919 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0.0029f
C4920 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.93e-21
C4921 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.54e-20
C4922 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 0.00106f
C4923 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# V_GND 0.0172f
C4924 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.0913f
C4925 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# V_GND 0.00592f
C4926 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00747f
C4927 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nor2_1_0/Y 0.018f
C4928 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# 4.42e-20
C4929 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__conb_1_42/HI -9.48e-19
C4930 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# -0.0594f
C4931 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# V_GND 0.00491f
C4932 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__nand2_8_9/Y 1.57e-19
C4933 sky130_fd_sc_hd__inv_1_18/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0138f
C4934 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_93/A 9.66e-20
C4935 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_27/LO 0.0474f
C4936 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# V_GND 1.67e-19
C4937 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00226f
C4938 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_581_47# -7.91e-19
C4939 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__inv_16_2/Y 0.00104f
C4940 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.08e-20
C4941 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.04e-21
C4942 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# V_LOW 1.62e-19
C4943 sky130_fd_sc_hd__conb_1_11/HI sky130_fd_sc_hd__inv_16_2/Y 0.0014f
C4944 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.578f
C4945 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_97/Y 0.00585f
C4946 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# sky130_fd_sc_hd__conb_1_27/HI 2e-19
C4947 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_17/Y 0.458f
C4948 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# sky130_fd_sc_hd__inv_1_60/Y 7.97e-21
C4949 sky130_fd_sc_hd__conb_1_26/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 5.51e-20
C4950 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# V_LOW -0.00266f
C4951 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# -0.00618f
C4952 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# V_LOW 0.0123f
C4953 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 2.89e-20
C4954 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 2.89e-20
C4955 sky130_fd_sc_hd__dfbbn_1_10/Q_N V_GND -0.00784f
C4956 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# sky130_fd_sc_hd__conb_1_9/HI -0.00125f
C4957 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__conb_1_36/HI 5.94e-19
C4958 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_16_2/Y 1.72e-20
C4959 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# V_LOW -0.0148f
C4960 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# V_LOW 0.0106f
C4961 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# sky130_fd_sc_hd__inv_1_22/Y 1.83e-20
C4962 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# V_GND 3.16e-19
C4963 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.24e-19
C4964 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 0.00304f
C4965 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_13/HI 2.23e-21
C4966 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# V_LOW 0.00334f
C4967 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# V_GND 0.00226f
C4968 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__inv_1_12/Y 0.00284f
C4969 sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# V_GND 1.77e-19
C4970 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_581_47# -2.6e-20
C4971 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# V_LOW 1.79e-20
C4972 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.64e-20
C4973 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# -0.00117f
C4974 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 4.48e-19
C4975 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# -9.88e-20
C4976 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# -0.00175f
C4977 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__conb_1_45/HI -2.17e-19
C4978 sky130_fd_sc_hd__nand2_8_3/Y V_LOW 0.245f
C4979 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 9.92e-21
C4980 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 4.44e-20
C4981 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 2.26e-21
C4982 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 1.51e-20
C4983 sky130_fd_sc_hd__dfbbn_1_12/a_581_47# V_GND -9.16e-19
C4984 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 6.04e-20
C4985 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_9/Y 0.00281f
C4986 sky130_fd_sc_hd__dfbbn_1_39/Q_N FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0237f
C4987 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_21/HI 2.56e-20
C4988 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# -4.66e-20
C4989 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# V_LOW 2.26e-20
C4990 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# -2.32e-19
C4991 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -0.00148f
C4992 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__conb_1_37/HI 1.1e-21
C4993 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 7.13e-21
C4994 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# V_GND 1.76e-19
C4995 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# V_GND -0.00195f
C4996 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_71/A 4.43e-21
C4997 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 0.0134f
C4998 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 9.74e-22
C4999 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 1.34e-20
C5000 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_1_99/Y 0.031f
C5001 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# 0.00306f
C5002 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_93/A 1.32e-19
C5003 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# V_GND -0.00614f
C5004 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# V_LOW 2.26e-20
C5005 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# V_LOW 4.8e-20
C5006 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__conb_1_44/HI 4.47e-20
C5007 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 0.013f
C5008 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# V_GND -3.81e-19
C5009 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_12/Y 2.91e-21
C5010 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# V_LOW -0.00266f
C5011 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.1e-21
C5012 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.64e-19
C5013 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# 1.48e-19
C5014 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# V_LOW -0.00149f
C5015 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# V_GND 0.00172f
C5016 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__conb_1_41/LO 1.12e-19
C5017 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_1/LO 0.00126f
C5018 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# Reset 0.00427f
C5019 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.04e-19
C5020 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# V_GND 0.00155f
C5021 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__conb_1_41/HI 3.27e-21
C5022 sky130_fd_sc_hd__conb_1_24/LO V_LOW 0.0971f
C5023 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/Q_N 0.0252f
C5024 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_8_6/a_27_47# 0.00103f
C5025 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_381_47# -0.00441f
C5026 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# Reset 0.00825f
C5027 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_16/HI 3.66e-20
C5028 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 5.74e-20
C5029 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 4.14e-21
C5030 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# V_GND -0.00444f
C5031 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.427f
C5032 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__inv_1_21/Y 2.46e-19
C5033 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# 0.00174f
C5034 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# V_GND 2.63e-19
C5035 sky130_fd_sc_hd__dfbbn_1_38/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 6.42e-19
C5036 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__conb_1_42/HI -2.17e-19
C5037 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# V_GND 2.41e-19
C5038 sky130_fd_sc_hd__conb_1_46/LO V_LOW 0.0394f
C5039 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_193_47# -0.032f
C5040 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0354f
C5041 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_101/Y 7.23e-20
C5042 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# V_LOW -0.00121f
C5043 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_97/A 0.00432f
C5044 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 0.00885f
C5045 RISING_COUNTER.COUNT_SUB_DFF12.Q V_LOW 0.179f
C5046 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__conb_1_25/LO 4.55e-20
C5047 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__inv_1_19/Y 4.43e-21
C5048 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# -0.117f
C5049 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0.00163f
C5050 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0.00949f
C5051 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 0.00163f
C5052 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 7.67e-19
C5053 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 7.67e-19
C5054 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 0.00949f
C5055 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00675f
C5056 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.91e-19
C5057 sky130_fd_sc_hd__inv_1_26/Y V_SENSE 0.0957f
C5058 sky130_fd_sc_hd__conb_1_35/LO V_LOW 0.0659f
C5059 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_581_47# -7.91e-19
C5060 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_647_21# -0.00108f
C5061 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.285f
C5062 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 8.46e-19
C5063 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.00109f
C5064 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.00109f
C5065 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 3.97e-19
C5066 sky130_fd_sc_hd__dfbbn_1_46/Q_N sky130_fd_sc_hd__conb_1_36/HI -2.17e-19
C5067 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__conb_1_44/HI 0.0121f
C5068 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 4.85e-21
C5069 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 2.78e-20
C5070 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# V_LOW -0.0034f
C5071 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# V_LOW 2.94e-20
C5072 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# V_GND 0.00188f
C5073 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00186f
C5074 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 3.8e-21
C5075 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 1.26e-19
C5076 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__inv_1_65/Y 0.0112f
C5077 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 5.41e-21
C5078 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 3.43e-21
C5079 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 7.84e-21
C5080 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_49/HI 1.47e-19
C5081 sky130_fd_sc_hd__dfbbn_1_48/Q_N V_GND -0.00115f
C5082 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.3e-20
C5083 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.11e-19
C5084 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_557_413# 8.26e-19
C5085 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# V_LOW -0.312f
C5086 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 0.497f
C5087 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__nand3_1_2/Y 0.106f
C5088 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.41e-20
C5089 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# V_LOW 1.38e-19
C5090 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_557_413# 7.19e-19
C5091 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_41/HI -0.00128f
C5092 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__conb_1_15/LO 0.0116f
C5093 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# -1.64e-19
C5094 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_1_76/A 0.00187f
C5095 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 3.21e-21
C5096 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# sky130_fd_sc_hd__conb_1_32/HI 5.21e-19
C5097 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.33e-19
C5098 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__conb_1_40/LO 1.82e-19
C5099 sky130_fd_sc_hd__inv_1_70/A sky130_fd_sc_hd__inv_1_65/Y 4.48e-20
C5100 sky130_fd_sc_hd__inv_1_68/A sky130_fd_sc_hd__nand2_8_9/Y 9.77e-19
C5101 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# V_LOW -0.00121f
C5102 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# V_GND -0.00124f
C5103 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0354f
C5104 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_74/Y 4.05e-19
C5105 sky130_fd_sc_hd__inv_1_16/Y V_GND 0.0824f
C5106 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 3.63e-21
C5107 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 1.65e-20
C5108 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 7.67e-19
C5109 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 5.98e-19
C5110 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 7e-19
C5111 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 8.23e-19
C5112 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 7.07e-19
C5113 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -3.48e-20
C5114 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_891_329# -2.2e-20
C5115 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__conb_1_15/LO 9.17e-19
C5116 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 8.48e-19
C5117 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# 3.32e-19
C5118 sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# sky130_fd_sc_hd__conb_1_44/HI -6.57e-19
C5119 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_67/Y 1.67e-20
C5120 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.3e-19
C5121 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# V_GND 0.0199f
C5122 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# V_GND 9.17e-19
C5123 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.25e-20
C5124 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__inv_1_57/Y 3.32e-20
C5125 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00193f
C5126 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# Reset 1.51e-20
C5127 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 5.97e-21
C5128 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.00115f
C5129 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00241f
C5130 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.00192f
C5131 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 4.4e-20
C5132 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 3.82e-20
C5133 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# V_GND -0.00336f
C5134 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 1.42e-20
C5135 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# 0.00366f
C5136 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# -0.00138f
C5137 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -5.54e-21
C5138 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# -0.00141f
C5139 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00457f
C5140 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 9.14e-19
C5141 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 7.34e-19
C5142 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 1e-19
C5143 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0549f
C5144 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00523f
C5145 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_75/A 4.05e-20
C5146 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# -4.1e-19
C5147 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_891_329# -2.2e-20
C5148 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# V_GND 9.33e-19
C5149 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__inv_1_12/Y 2.35e-21
C5150 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__conb_1_51/HI 0.00321f
C5151 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0397f
C5152 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_95/A 3.29e-20
C5153 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 6e-19
C5154 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_76/A 0.00599f
C5155 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 4.85e-21
C5156 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 1.44e-19
C5157 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 0.036f
C5158 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_105/Y 0.0266f
C5159 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 0.00293f
C5160 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_1_12/Y 4.91e-19
C5161 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 8.18e-19
C5162 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 1.79e-19
C5163 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 1.99e-19
C5164 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_581_47# -2.6e-20
C5165 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00274f
C5166 sky130_fd_sc_hd__inv_1_58/Y sky130_fd_sc_hd__conb_1_26/HI 0.00238f
C5167 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# V_LOW -0.00526f
C5168 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0989f
C5169 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# -6.43e-20
C5170 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# -0.0133f
C5171 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 0.00127f
C5172 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# V_LOW 0.0183f
C5173 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# CLOCK_GEN.SR_Op.Q 4.88e-21
C5174 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_1_112/Y 6.56e-19
C5175 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__conb_1_36/HI 2.06e-20
C5176 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 2.59e-19
C5177 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.0732f
C5178 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF9.Q 1.33f
C5179 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__inv_16_0/Y 8.65e-19
C5180 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# V_LOW 0.0148f
C5181 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0106f
C5182 Reset sky130_fd_sc_hd__inv_1_68/A 1.47e-20
C5183 transmission_gate_0/GN sky130_fd_sc_hd__inv_2_0/Y 0.214f
C5184 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 6.82e-20
C5185 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# V_GND 0.00627f
C5186 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 1.16e-19
C5187 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__conb_1_40/HI 1.44e-21
C5188 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 0.0239f
C5189 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.78e-22
C5190 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 5.41e-21
C5191 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 8.79e-22
C5192 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__inv_1_53/Y 2.96e-20
C5193 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__inv_1_13/Y 3.95e-19
C5194 sky130_fd_sc_hd__inv_1_85/Y Reset 0.167f
C5195 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_70/Y 0.00228f
C5196 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# V_GND -0.00474f
C5197 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__conb_1_41/HI -4.01e-20
C5198 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 0.00319f
C5199 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 0.00166f
C5200 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__conb_1_13/LO 1.88e-19
C5201 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# V_GND 0.00421f
C5202 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.075f
C5203 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 2.26e-19
C5204 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 0.00106f
C5205 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 2.26e-19
C5206 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0.00803f
C5207 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0.00106f
C5208 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_18/LO 5.28e-21
C5209 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# V_GND 0.00495f
C5210 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 3.48e-20
C5211 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# -0.00142f
C5212 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00163f
C5213 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 7.8e-21
C5214 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__inv_1_103/Y 0.0173f
C5215 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_47/HI 0.336f
C5216 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# V_GND 4.98e-19
C5217 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_1_108/Y 5.16e-19
C5218 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_16_0/Y 2.5e-20
C5219 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__conb_1_27/HI 1.14e-20
C5220 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_891_329# -0.0016f
C5221 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# -0.00492f
C5222 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# V_LOW 4.8e-20
C5223 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.68e-20
C5224 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 5.03e-19
C5225 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 9.74e-19
C5226 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__conb_1_40/HI 0.0268f
C5227 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 0.00491f
C5228 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 3.66e-20
C5229 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_1_54/Y 1.9e-20
C5230 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_85/A 0.45f
C5231 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 1.07e-21
C5232 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 5.73e-20
C5233 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# -9.32e-20
C5234 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.9e-19
C5235 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 5.21e-19
C5236 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# sky130_fd_sc_hd__inv_16_1/Y 2.45e-19
C5237 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0548f
C5238 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__inv_1_23/Y 0.00667f
C5239 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_16_0/Y 0.309f
C5240 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_1_90/Y 5.81e-20
C5241 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_76/A 4.38e-19
C5242 sky130_fd_sc_hd__inv_1_100/Y sky130_fd_sc_hd__inv_16_1/Y 0.0225f
C5243 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_9/Y 2.55e-20
C5244 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 7.13e-20
C5245 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__inv_1_98/Y 9.48e-20
C5246 sky130_fd_sc_hd__dfbbn_1_49/a_581_47# V_GND 2.24e-19
C5247 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 7.76e-20
C5248 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# sky130_fd_sc_hd__conb_1_51/HI 3.95e-21
C5249 sky130_fd_sc_hd__dfbbn_1_7/Q_N FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0143f
C5250 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# 4.48e-21
C5251 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 7.06e-19
C5252 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 5.4e-20
C5253 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 3.2e-21
C5254 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 8.88e-19
C5255 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 5.15e-19
C5256 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 4.94e-20
C5257 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.00596f
C5258 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 6.4e-19
C5259 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__inv_1_54/Y 2.48e-20
C5260 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# V_LOW 4.8e-20
C5261 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 8.65e-20
C5262 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_581_47# 1.4e-19
C5263 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 7.3e-19
C5264 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# 6.06e-21
C5265 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 1.1e-20
C5266 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_33/LO 1.85e-21
C5267 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.0474f
C5268 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/Q_N 1.76e-19
C5269 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 1.76e-19
C5270 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__conb_1_23/HI 1.88e-19
C5271 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 4.56e-21
C5272 FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_35/HI 0.0258f
C5273 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.166f
C5274 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.00101f
C5275 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 5.8e-19
C5276 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 2.11e-19
C5277 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_791_47# 5.72e-20
C5278 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 1.79e-20
C5279 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 6.34e-20
C5280 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 4.55e-20
C5281 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 4.49e-21
C5282 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 7.33e-20
C5283 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00128f
C5284 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 3.55e-20
C5285 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__conb_1_46/HI -0.0139f
C5286 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__conb_1_2/HI 0.00399f
C5287 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.554f
C5288 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00116f
C5289 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__inv_1_103/Y 0.0144f
C5290 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# V_LOW 2.94e-20
C5291 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_100/Y 4.91e-19
C5292 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 4.85e-21
C5293 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.00478f
C5294 sky130_fd_sc_hd__dfbbn_1_17/a_581_47# V_GND 2.41e-19
C5295 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.51e-20
C5296 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_8/LO 0.00268f
C5297 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# 0.0169f
C5298 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 2.81e-20
C5299 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 1.38e-19
C5300 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 0.00478f
C5301 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.00256f
C5302 sky130_fd_sc_hd__conb_1_33/HI V_GND 0.164f
C5303 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 4.68e-21
C5304 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00645f
C5305 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# V_LOW 0.0608f
C5306 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# sky130_fd_sc_hd__inv_1_53/Y 3.37e-19
C5307 FULL_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 2.06e-19
C5308 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# V_GND -0.00511f
C5309 sky130_fd_sc_hd__inv_1_80/A V_GND 0.348f
C5310 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 2.65e-22
C5311 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 5.11e-20
C5312 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 5.03e-20
C5313 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 6.48e-20
C5314 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_791_47# 8.71e-19
C5315 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_40/A 0.0443f
C5316 sky130_fd_sc_hd__nand2_8_0/a_27_47# V_LOW -0.00471f
C5317 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 3.55e-19
C5318 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__inv_1_17/Y 7.61e-20
C5319 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# V_GND 6.86e-19
C5320 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# -5.54e-21
C5321 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -2.6e-19
C5322 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# -3.8e-20
C5323 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.045f
C5324 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_473_413# 2.68e-20
C5325 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# 1.5e-19
C5326 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 1.5e-19
C5327 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# V_GND 0.00156f
C5328 sky130_fd_sc_hd__nand3_1_2/B sky130_fd_sc_hd__inv_1_75/A 0.0257f
C5329 sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__nand2_8_2/A 3.85e-20
C5330 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# 9.28e-19
C5331 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 3.4e-20
C5332 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 3.61e-20
C5333 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 3.4e-20
C5334 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 7.07e-20
C5335 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# sky130_fd_sc_hd__conb_1_27/HI 5.52e-20
C5336 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# -0.00282f
C5337 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# V_GND 0.00396f
C5338 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_891_329# -0.00159f
C5339 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# -0.00279f
C5340 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_47/Y 2.55e-21
C5341 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 1.36e-19
C5342 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00399f
C5343 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# sky130_fd_sc_hd__conb_1_35/HI 5.75e-19
C5344 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# Reset 1.75e-19
C5345 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.00184f
C5346 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_23/Y 2.04e-22
C5347 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# sky130_fd_sc_hd__conb_1_45/HI 7.28e-19
C5348 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.37e-19
C5349 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/Q_N -4.33e-20
C5350 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 4.15e-19
C5351 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.99e-20
C5352 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 4.4e-19
C5353 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 4.78e-20
C5354 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_107/Y 4.94e-21
C5355 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_39/LO 3.05e-20
C5356 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00359f
C5357 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.06e-20
C5358 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_93/Y 0.00236f
C5359 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__conb_1_0/HI 3.27e-19
C5360 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__nand2_1_5/a_113_47# 7.29e-19
C5361 sky130_fd_sc_hd__conb_1_44/LO sky130_fd_sc_hd__conb_1_44/HI 0.00337f
C5362 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0144f
C5363 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_193_47# 2.51e-20
C5364 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.3e-20
C5365 sky130_fd_sc_hd__inv_1_56/Y sky130_fd_sc_hd__inv_1_57/Y 4.73e-21
C5366 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00613f
C5367 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 2.18e-20
C5368 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.37e-20
C5369 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 9.94e-20
C5370 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_16_0/Y 4.38e-19
C5371 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 0.00137f
C5372 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/Q_N 0.026f
C5373 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.0638f
C5374 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 1.81e-20
C5375 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 1.29e-19
C5376 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00237f
C5377 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 4.97e-19
C5378 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.00105f
C5379 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_17/HI 0.0213f
C5380 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 7.24e-21
C5381 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__nand2_8_2/A 0.072f
C5382 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 8.93e-20
C5383 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__conb_1_33/HI -5.12e-20
C5384 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# sky130_fd_sc_hd__conb_1_2/HI -1.17e-19
C5385 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# -5.54e-21
C5386 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__nand3_1_1/Y 3.99e-20
C5387 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# sky130_fd_sc_hd__inv_1_103/Y 6.02e-19
C5388 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_95/A 0.0765f
C5389 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_96/Y 0.0184f
C5390 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_20/Y 0.0709f
C5391 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 8.16e-19
C5392 RISING_COUNTER.COUNT_SUB_DFF10.Q V_GND 2.51f
C5393 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 9.03e-21
C5394 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 9.7e-20
C5395 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# 8.18e-21
C5396 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_78/A 4.43e-21
C5397 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 8.11e-21
C5398 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__conb_1_21/HI 5.31e-20
C5399 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0183f
C5400 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 0.00112f
C5401 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# V_LOW 1.61e-19
C5402 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# V_LOW -0.00576f
C5403 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 6.21e-21
C5404 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# V_LOW 2.94e-20
C5405 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# V_LOW 0.0244f
C5406 sky130_fd_sc_hd__dfbbn_1_5/Q_N V_GND -0.00751f
C5407 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 5.58e-21
C5408 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_941_21# -0.00147f
C5409 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# -2.28e-19
C5410 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_100/Y -7.56e-19
C5411 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0155f
C5412 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 0.014f
C5413 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# V_LOW -0.00376f
C5414 sky130_fd_sc_hd__conb_1_22/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 4.97e-20
C5415 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 1.51e-19
C5416 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# 4.82e-19
C5417 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# -9.32e-20
C5418 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_68/Y 1.02e-20
C5419 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0265f
C5420 FALLING_COUNTER.COUNT_SUB_DFF10.Q V_GND 0.999f
C5421 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_381_47# 4.39e-19
C5422 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 4.39e-19
C5423 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# V_LOW 1.38e-19
C5424 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# V_GND 5.08e-19
C5425 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# V_GND 1.4e-19
C5426 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# V_LOW 0.0153f
C5427 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__conb_1_27/HI 6.55e-19
C5428 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__conb_1_28/LO 6.23e-21
C5429 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_381_47# -2.53e-20
C5430 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_557_413# 0.00216f
C5431 sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# V_GND 4.62e-19
C5432 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# V_GND 2.42e-19
C5433 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# -0.00385f
C5434 sky130_fd_sc_hd__nand2_1_1/a_113_47# V_LOW -1.78e-19
C5435 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_37/LO 1.79e-19
C5436 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_106/Y 0.182f
C5437 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# V_GND 5.83e-19
C5438 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_473_413# -0.012f
C5439 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -0.00932f
C5440 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# V_LOW 0.049f
C5441 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.00326f
C5442 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.015f
C5443 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00252f
C5444 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 2.3e-19
C5445 sky130_fd_sc_hd__dfbbn_1_47/Q_N RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0225f
C5446 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -0.00932f
C5447 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_473_413# -0.0127f
C5448 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# 8.95e-21
C5449 FULL_COUNTER.COUNT_SUB_DFF16.Q V_GND 1.68f
C5450 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_1/Y 0.37f
C5451 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__conb_1_49/HI 4.12e-21
C5452 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF1.Q 3.66e-20
C5453 sky130_fd_sc_hd__conb_1_10/LO FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0143f
C5454 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 5.32e-20
C5455 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# V_GND 7.65e-19
C5456 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 5.1e-21
C5457 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_1_59/Y 4.49e-19
C5458 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0827f
C5459 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# V_GND 0.00188f
C5460 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# Reset 0.00137f
C5461 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.89e-19
C5462 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.14e-20
C5463 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0321f
C5464 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__inv_1_61/Y 1.44e-19
C5465 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00115f
C5466 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_32/A 1.98e-20
C5467 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_32/Y 4.38e-19
C5468 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# V_LOW 1.38e-19
C5469 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# V_GND 0.00413f
C5470 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/Q_N 5.88e-21
C5471 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 0.00193f
C5472 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# -0.148f
C5473 sky130_fd_sc_hd__inv_1_45/Y V_LOW 0.0925f
C5474 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00379f
C5475 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__conb_1_41/HI 2.23e-20
C5476 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00202f
C5477 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__inv_1_4/Y 0.00227f
C5478 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/Q_N 1.15e-19
C5479 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.51e-21
C5480 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__conb_1_33/HI -2.07e-19
C5481 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.15e-20
C5482 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.22e-20
C5483 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# Reset 2.68e-19
C5484 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00789f
C5485 sky130_fd_sc_hd__conb_1_4/LO V_GND 0.00933f
C5486 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# -2.35e-19
C5487 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -1.89e-19
C5488 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# sky130_fd_sc_hd__inv_16_2/Y 2.57e-20
C5489 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 8.86e-21
C5490 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 7.45e-21
C5491 sky130_fd_sc_hd__conb_1_32/HI V_GND -0.141f
C5492 sky130_fd_sc_hd__nand2_8_3/Y sky130_fd_sc_hd__inv_1_80/A 0.00426f
C5493 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_21/LO 0.00297f
C5494 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# -0.0213f
C5495 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_557_413# -0.0012f
C5496 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__inv_1_58/Y 9.77e-20
C5497 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# V_GND 8.42e-19
C5498 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# sky130_fd_sc_hd__inv_1_11/Y 1.96e-20
C5499 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.21e-21
C5500 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/Q_N 4.43e-20
C5501 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 2.25e-20
C5502 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.49e-21
C5503 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# V_LOW 0.00586f
C5504 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_75/A 0.00508f
C5505 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__conb_1_8/HI 0.00148f
C5506 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# V_LOW 0.0114f
C5507 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# -7.17e-20
C5508 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# -1.64e-19
C5509 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.00103f
C5510 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 7.29e-19
C5511 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# V_LOW 0.0113f
C5512 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 5.62e-19
C5513 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_24/HI 5.95e-21
C5514 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/Q_N -4.78e-20
C5515 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__conb_1_13/HI 6.53e-19
C5516 sky130_fd_sc_hd__inv_1_55/Y V_LOW 0.23f
C5517 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0101f
C5518 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00524f
C5519 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_25/HI 0.0263f
C5520 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 8.84e-20
C5521 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0361f
C5522 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00148f
C5523 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__inv_1_17/Y 0.00773f
C5524 sky130_fd_sc_hd__dfbbn_1_44/a_1672_329# V_LOW 1.79e-20
C5525 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__inv_1_105/Y 0.0174f
C5526 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# -1.44e-20
C5527 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00648f
C5528 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# V_GND 0.00183f
C5529 sky130_fd_sc_hd__conb_1_50/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 2.48e-20
C5530 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_21/HI 3.27e-19
C5531 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/Q_N -4.97e-19
C5532 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# sky130_fd_sc_hd__conb_1_28/HI 8.98e-20
C5533 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# -0.0494f
C5534 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# V_LOW 2.94e-20
C5535 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.3e-19
C5536 sky130_fd_sc_hd__dfbbn_1_19/a_557_413# V_GND 1.72e-19
C5537 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# -2.57e-20
C5538 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# CLOCK_GEN.SR_Op.Q 1.33e-19
C5539 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 4.73e-19
C5540 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.0427f
C5541 sky130_fd_sc_hd__fill_4_56/VPB V_LOW 0.797f
C5542 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 5.88e-19
C5543 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 7.67e-19
C5544 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0.00863f
C5545 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 8.42e-19
C5546 sky130_fd_sc_hd__inv_1_100/Y V_LOW 0.217f
C5547 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.58e-19
C5548 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# -2.57e-20
C5549 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_647_21# -0.00115f
C5550 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 6.57e-20
C5551 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__conb_1_39/LO 2.14e-19
C5552 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.00119f
C5553 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_72/A 6.97e-20
C5554 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.76e-21
C5555 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# sky130_fd_sc_hd__conb_1_49/HI -2.65e-20
C5556 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.87e-20
C5557 Reset V_HIGH 0.186f
C5558 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__inv_1_59/Y 3.75e-20
C5559 sky130_fd_sc_hd__dfbbn_1_44/a_1363_47# V_GND 1.88e-19
C5560 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# 8.66e-21
C5561 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# Reset 4.54e-19
C5562 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 1.25e-19
C5563 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00122f
C5564 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__inv_1_61/Y 3.01e-19
C5565 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00225f
C5566 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 3.62e-21
C5567 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# 9.06e-20
C5568 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# V_GND 0.0273f
C5569 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.014f
C5570 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_557_413# -0.0012f
C5571 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# -0.0105f
C5572 sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF10.Q 9.87e-20
C5573 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# V_GND 6.11e-19
C5574 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.402f
C5575 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_67/Y 2.15e-20
C5576 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__inv_16_2/Y 0.428f
C5577 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_20/HI 4.37e-19
C5578 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_0/Y 0.484f
C5579 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 4.04e-20
C5580 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.00379f
C5581 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 8.74e-19
C5582 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 0.00208f
C5583 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0.00208f
C5584 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 3.53e-19
C5585 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/Q_N -4.78e-20
C5586 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.22e-21
C5587 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_94/A 0.00131f
C5588 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# -6.43e-20
C5589 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# -3.06e-20
C5590 sky130_fd_sc_hd__inv_1_52/Y CLOCK_GEN.SR_Op.Q 3.68e-19
C5591 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 7.69e-20
C5592 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 1.5e-19
C5593 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# -1.66e-19
C5594 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.00386f
C5595 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 1.04e-19
C5596 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# -6.23e-21
C5597 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# -0.00527f
C5598 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_10/Y 0.00819f
C5599 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# -5.42e-19
C5600 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# sky130_fd_sc_hd__inv_1_60/Y 5.15e-21
C5601 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.91e-19
C5602 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 3.19e-19
C5603 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.029f
C5604 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# -0.0309f
C5605 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_557_413# -3.67e-20
C5606 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF1.Q 4.5e-19
C5607 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/Q_N 0.00482f
C5608 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 8.5e-21
C5609 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__conb_1_8/HI 4.4e-19
C5610 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 0.00472f
C5611 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# V_LOW -0.00121f
C5612 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_557_413# -0.0012f
C5613 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_891_329# -1.42e-19
C5614 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# -0.00393f
C5615 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00184f
C5616 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0156f
C5617 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 7.1e-19
C5618 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_105/Y 0.035f
C5619 sky130_fd_sc_hd__inv_1_103/Y sky130_fd_sc_hd__conb_1_45/HI 0.00544f
C5620 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_43/A 0.0461f
C5621 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.00144f
C5622 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 1.9e-20
C5623 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# V_LOW 0.0043f
C5624 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_28/HI 5.61e-19
C5625 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__inv_1_15/Y 7.53e-19
C5626 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.01e-20
C5627 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__inv_1_5/Y 0.00592f
C5628 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__conb_1_13/HI 0.00128f
C5629 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_103/Y 0.0479f
C5630 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 6.15e-21
C5631 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 3.9e-21
C5632 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 2.63e-21
C5633 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.37e-19
C5634 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 3.22e-21
C5635 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 3.97e-22
C5636 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.05e-21
C5637 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_2/LO 0.00366f
C5638 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__inv_1_90/Y 1.07e-20
C5639 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 8.78e-20
C5640 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# sky130_fd_sc_hd__conb_1_25/HI 3.6e-19
C5641 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__inv_1_9/Y 0.00198f
C5642 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.35e-20
C5643 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.71e-21
C5644 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.159f
C5645 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# V_GND 0.00167f
C5646 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.237f
C5647 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 0.00144f
C5648 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# V_LOW 2.26e-20
C5649 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__conb_1_37/HI -1.14e-20
C5650 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.45e-19
C5651 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# 7.08e-20
C5652 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 0.00488f
C5653 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 9.28e-20
C5654 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.274f
C5655 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.48e-19
C5656 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 3.1e-19
C5657 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 0.00243f
C5658 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.3e-19
C5659 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 1.6e-21
C5660 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 1.48e-22
C5661 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 5.43e-20
C5662 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_581_47# -7.91e-19
C5663 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_1/a_381_47# 8.6e-20
C5664 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 8.68e-20
C5665 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.03e-20
C5666 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# sky130_fd_sc_hd__inv_1_19/Y 0.00147f
C5667 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# 4.03e-19
C5668 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 4.84e-20
C5669 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_48/LO 6.98e-21
C5670 sky130_fd_sc_hd__conb_1_46/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0278f
C5671 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 2.68e-21
C5672 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# V_GND 0.00213f
C5673 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__conb_1_19/HI 0.0649f
C5674 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__conb_1_28/LO 1.03e-19
C5675 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_97/Y 1.6e-19
C5676 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__conb_1_6/HI 2.67e-19
C5677 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# sky130_fd_sc_hd__conb_1_20/HI 0.00557f
C5678 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 4.43e-21
C5679 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_6/HI 0.0373f
C5680 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 3.63e-19
C5681 sky130_fd_sc_hd__conb_1_18/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0106f
C5682 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 9.65e-19
C5683 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 7.56e-20
C5684 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0.00111f
C5685 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 1.34e-20
C5686 sky130_fd_sc_hd__inv_1_99/Y V_GND 0.136f
C5687 sky130_fd_sc_hd__dfbbn_1_28/Q_N RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0294f
C5688 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# -6.57e-19
C5689 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 0.00114f
C5690 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_95/Y 2.95e-19
C5691 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_18/Y 0.0313f
C5692 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_41/LO 6.46e-20
C5693 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 6.27e-20
C5694 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# 0.0023f
C5695 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 1.44e-19
C5696 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 2.7e-20
C5697 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 5.52e-19
C5698 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00803f
C5699 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.00116f
C5700 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 6.94e-19
C5701 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.11e-20
C5702 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 0.00222f
C5703 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_17/HI 3.9e-20
C5704 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 4.09e-20
C5705 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# V_LOW -0.00389f
C5706 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__inv_1_53/Y 8.84e-19
C5707 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.25e-20
C5708 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0679f
C5709 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 0.00412f
C5710 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__conb_1_11/HI 5.52e-20
C5711 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.141f
C5712 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__conb_1_8/HI 5.86e-19
C5713 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand3_1_0/Y 0.33f
C5714 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.131f
C5715 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0329f
C5716 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# CLOCK_GEN.SR_Op.Q 2.46e-20
C5717 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00959f
C5718 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__inv_1_15/Y 1.28e-20
C5719 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 7.3e-22
C5720 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# CLOCK_GEN.SR_Op.Q 0.0293f
C5721 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# V_LOW -2.54e-19
C5722 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 4.52e-21
C5723 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0291f
C5724 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 2.89e-21
C5725 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 5.55e-19
C5726 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0158f
C5727 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__conb_1_12/HI 6.26e-21
C5728 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# V_GND 7.65e-19
C5729 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 7.23e-19
C5730 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1_21/HI 4.17e-19
C5731 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 0.00704f
C5732 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00304f
C5733 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 1.46e-20
C5734 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 3.45e-20
C5735 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__conb_1_31/HI 2.61e-19
C5736 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__conb_1_31/HI 7.75e-21
C5737 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__conb_1_26/HI 1.62e-19
C5738 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# sky130_fd_sc_hd__conb_1_37/HI -3.05e-20
C5739 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 1.75e-20
C5740 FALLING_COUNTER.COUNT_SUB_DFF2.Q V_LOW 2.09f
C5741 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.31e-20
C5742 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 0.00117f
C5743 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 7.45e-21
C5744 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 2.55e-19
C5745 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0136f
C5746 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# 0.00165f
C5747 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.16e-20
C5748 sky130_fd_sc_hd__conb_1_34/LO V_GND 0.00108f
C5749 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_75/A 7.14e-20
C5750 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 8.74e-21
C5751 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# V_GND 0.0121f
C5752 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 1.94e-20
C5753 sky130_fd_sc_hd__dfbbn_1_40/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.13e-20
C5754 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_112/Y 1.82e-20
C5755 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__inv_16_1/Y 0.442f
C5756 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_64/A 0.115f
C5757 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 0.00141f
C5758 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__conb_1_42/HI 6.75e-19
C5759 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_51/LO 0.00371f
C5760 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_8/Y 0.00656f
C5761 sky130_fd_sc_hd__inv_1_75/A sky130_fd_sc_hd__nand2_8_2/A 0.087f
C5762 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_93/Y 0.00183f
C5763 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# sky130_fd_sc_hd__conb_1_5/HI 4.7e-20
C5764 sky130_fd_sc_hd__conb_1_45/LO V_GND -0.00454f
C5765 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_47/Y 0.00532f
C5766 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 0.032f
C5767 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__conb_1_21/LO 1.38e-21
C5768 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__conb_1_21/HI 0.00395f
C5769 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 8.79e-20
C5770 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 7.26e-19
C5771 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_16/HI 1.65e-19
C5772 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.00102f
C5773 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0.00145f
C5774 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_647_21# -1.24e-20
C5775 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_1_9/Y 5.09e-20
C5776 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_66/Y 0.0069f
C5777 sky130_fd_sc_hd__conb_1_43/HI V_GND 0.309f
C5778 sky130_fd_sc_hd__inv_1_34/A V_GND 0.0807f
C5779 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 1.3e-21
C5780 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_22/Y 4.43e-21
C5781 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_98/Y 0.337f
C5782 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 3.35e-19
C5783 sky130_fd_sc_hd__dfbbn_1_44/Q_N RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00266f
C5784 sky130_fd_sc_hd__inv_1_94/Y V_GND 0.157f
C5785 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_29/LO 2.09e-20
C5786 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__inv_1_58/Y 4.27e-20
C5787 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 9.04e-20
C5788 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.051f
C5789 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00565f
C5790 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 3.79e-21
C5791 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 7.56e-20
C5792 sky130_fd_sc_hd__inv_1_56/Y RISING_COUNTER.COUNT_SUB_DFF15.Q 1.13e-19
C5793 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_112/Y 0.222f
C5794 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.06e-21
C5795 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__conb_1_25/HI 9.44e-19
C5796 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.8e-19
C5797 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__conb_1_2/HI 2.27e-20
C5798 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.13e-21
C5799 RISING_COUNTER.COUNT_SUB_DFF8.Q V_GND 0.948f
C5800 sky130_fd_sc_hd__conb_1_0/HI V_GND 0.0399f
C5801 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__inv_1_101/Y 0.0167f
C5802 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 0.548f
C5803 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__inv_1_11/Y 1.75e-19
C5804 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__conb_1_30/HI 3.26e-20
C5805 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# -6.43e-20
C5806 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# -3.06e-20
C5807 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0169f
C5808 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 4.26e-21
C5809 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.11e-20
C5810 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 7.72e-22
C5811 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 2.12e-21
C5812 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_1_90/Y 5.85e-22
C5813 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# 4.49e-21
C5814 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.00139f
C5815 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00244f
C5816 sky130_fd_sc_hd__dfbbn_1_28/a_557_413# sky130_fd_sc_hd__inv_1_54/Y 5.11e-19
C5817 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_13/LO 4.66e-21
C5818 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.22e-20
C5819 sky130_fd_sc_hd__nand3_1_2/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00503f
C5820 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__conb_1_39/HI 0.00378f
C5821 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 3.29e-19
C5822 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.0124f
C5823 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.00799f
C5824 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 6.02e-19
C5825 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00245f
C5826 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# V_LOW 0.00496f
C5827 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00987f
C5828 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__inv_1_11/Y 1.38e-19
C5829 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_791_47# 4.16e-20
C5830 sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# sky130_fd_sc_hd__conb_1_26/HI 0.00161f
C5831 sky130_fd_sc_hd__inv_1_18/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 2.88e-20
C5832 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_14/HI 0.0966f
C5833 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 5.06e-21
C5834 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.71e-19
C5835 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 0.0203f
C5836 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__inv_16_0/Y -3.75e-20
C5837 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 5.34e-20
C5838 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# 1.35e-20
C5839 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 4.54e-20
C5840 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# 2.42e-22
C5841 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00177f
C5842 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# -0.009f
C5843 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# V_GND 0.0086f
C5844 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.79e-19
C5845 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.464f
C5846 sky130_fd_sc_hd__conb_1_50/HI RISING_COUNTER.COUNT_SUB_DFF7.Q 1.55e-19
C5847 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00626f
C5848 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 0.016f
C5849 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 1.03e-19
C5850 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# CLOCK_GEN.SR_Op.Q 4.45e-20
C5851 sky130_fd_sc_hd__inv_1_119/Y V_LOW 0.601f
C5852 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__conb_1_22/HI 8.72e-19
C5853 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# V_LOW 0.00477f
C5854 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__conb_1_49/HI 2.67e-20
C5855 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_791_47# 5.96e-19
C5856 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# V_GND 0.01f
C5857 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_22/Y 1.33e-20
C5858 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0223f
C5859 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# V_LOW 0.0157f
C5860 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.21e-19
C5861 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 1.65e-19
C5862 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# V_LOW 0.0183f
C5863 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_37/LO 7.32e-21
C5864 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# V_GND -5.48e-19
C5865 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.72e-20
C5866 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__nand3_1_1/Y 0.118f
C5867 sky130_fd_sc_hd__inv_1_89/Y Reset 0.00424f
C5868 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_75/Y 0.00279f
C5869 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.86e-21
C5870 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 2.61e-20
C5871 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_557_413# -0.0012f
C5872 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_891_329# -2.46e-19
C5873 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# -0.0268f
C5874 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_581_47# -2.6e-20
C5875 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_1_6/Y 1.72e-20
C5876 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_1_107/Y 8.38e-20
C5877 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0139f
C5878 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.11e-21
C5879 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 9.65e-19
C5880 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__conb_1_18/HI 8.35e-20
C5881 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__inv_16_1/Y 0.0257f
C5882 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# V_GND 0.00719f
C5883 sky130_fd_sc_hd__conb_1_30/HI RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00202f
C5884 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# V_GND -0.0197f
C5885 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__conb_1_17/HI 8.03e-21
C5886 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0222f
C5887 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0.0127f
C5888 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__conb_1_23/HI -6.57e-19
C5889 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.64e-20
C5890 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# V_GND 0.00772f
C5891 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.63e-20
C5892 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_557_413# 4.16e-19
C5893 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__conb_1_28/HI -0.00218f
C5894 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_31/Y 0.0443f
C5895 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_2/Y 0.32f
C5896 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# sky130_fd_sc_hd__conb_1_25/HI -6.57e-19
C5897 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_11/HI 2.55e-20
C5898 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__inv_1_106/Y -3.15e-20
C5899 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# -5.54e-21
C5900 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# -0.00156f
C5901 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_16/HI 3.39e-19
C5902 sky130_fd_sc_hd__inv_1_14/Y V_LOW 0.0193f
C5903 sky130_fd_sc_hd__conb_1_6/LO V_GND -0.00531f
C5904 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# sky130_fd_sc_hd__conb_1_30/HI -0.00746f
C5905 sky130_fd_sc_hd__conb_1_23/HI CLOCK_GEN.SR_Op.Q 1.01e-20
C5906 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 2.37e-20
C5907 sky130_fd_sc_hd__inv_1_54/Y V_GND 0.013f
C5908 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_647_21# -0.00392f
C5909 sky130_fd_sc_hd__dfbbn_1_20/Q_N RISING_COUNTER.COUNT_SUB_DFF2.Q 9.19e-20
C5910 sky130_fd_sc_hd__conb_1_25/HI CLOCK_GEN.SR_Op.Q 0.0264f
C5911 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# V_LOW -0.0153f
C5912 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_381_47# 0.0109f
C5913 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__conb_1_10/HI 5.94e-19
C5914 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 0.00106f
C5915 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 5.77e-19
C5916 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# V_GND 0.00105f
C5917 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 4.23e-19
C5918 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# sky130_fd_sc_hd__conb_1_22/HI 4.09e-19
C5919 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF17.Q 0.0155f
C5920 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# V_GND -9.92e-20
C5921 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_15/Y 4.43e-21
C5922 FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_16_2/Y 0.27f
C5923 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -2.18e-19
C5924 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# -0.00263f
C5925 sky130_fd_sc_hd__dfbbn_1_2/a_581_47# sky130_fd_sc_hd__inv_1_76/A 1.58e-20
C5926 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# 3.59e-19
C5927 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__conb_1_16/HI 1.57e-20
C5928 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_1_18/Y 4.8e-19
C5929 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__conb_1_39/HI 6.77e-20
C5930 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00114f
C5931 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__inv_1_99/Y 8.73e-19
C5932 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# V_LOW 1.38e-19
C5933 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_381_47# 0.0107f
C5934 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__conb_1_12/HI 1.05e-19
C5935 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 1.34e-19
C5936 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# 3.22e-19
C5937 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# V_LOW -0.00121f
C5938 sky130_fd_sc_hd__conb_1_22/LO V_LOW 0.0949f
C5939 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.34e-19
C5940 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_581_47# -2.6e-20
C5941 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/Q_N 7.1e-20
C5942 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# V_GND -0.00279f
C5943 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.44e-19
C5944 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.89e-20
C5945 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 8.97e-20
C5946 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__conb_1_39/HI 0.00193f
C5947 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00201f
C5948 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# CLOCK_GEN.SR_Op.Q 2.47e-19
C5949 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_1_12/Y 5.9e-19
C5950 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# 2.82e-19
C5951 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 3.34e-19
C5952 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 3.74e-19
C5953 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__inv_1_18/Y 0.0304f
C5954 RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00111f
C5955 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# sky130_fd_sc_hd__conb_1_22/HI 4.61e-22
C5956 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.1e-20
C5957 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 7.01e-19
C5958 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# -3.51e-19
C5959 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# sky130_fd_sc_hd__inv_1_57/Y 9.74e-19
C5960 sky130_fd_sc_hd__conb_1_18/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00856f
C5961 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# V_GND 0.0108f
C5962 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# V_GND 7.97e-19
C5963 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0375f
C5964 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__inv_1_99/Y 0.00948f
C5965 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_45/HI 0.401f
C5966 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0012f
C5967 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_35/HI 0.0221f
C5968 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# V_GND 0.00312f
C5969 sky130_fd_sc_hd__conb_1_9/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 7.01e-21
C5970 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.22e-19
C5971 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 2.96e-19
C5972 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__inv_16_0/Y 9.99e-20
C5973 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# sky130_fd_sc_hd__conb_1_40/HI 0.00134f
C5974 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 4.81e-20
C5975 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 7.04e-19
C5976 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.0116f
C5977 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_71/A 0.0201f
C5978 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0285f
C5979 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 1.39e-19
C5980 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0193f
C5981 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__inv_16_1/Y 0.0413f
C5982 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0595f
C5983 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.15e-20
C5984 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__conb_1_44/HI 4.55e-21
C5985 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.5e-21
C5986 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# V_GND 0.00307f
C5987 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00795f
C5988 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__nand3_1_0/Y 7.07e-21
C5989 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__conb_1_18/HI -2.65e-20
C5990 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 1.83e-20
C5991 RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_28/HI 5.16e-20
C5992 sky130_fd_sc_hd__nand2_8_9/Y sky130_fd_sc_hd__inv_1_63/Y 0.0454f
C5993 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# V_GND 1.88e-19
C5994 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# V_LOW 2.26e-20
C5995 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__conb_1_17/HI 0.00149f
C5996 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__conb_1_38/HI 8.5e-21
C5997 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__inv_16_2/Y 8.53e-19
C5998 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# V_GND 3.04e-19
C5999 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 6.38e-21
C6000 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__nand3_1_0/Y 3.68e-19
C6001 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# V_LOW -0.00121f
C6002 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_473_413# 0.00978f
C6003 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__conb_1_45/HI 0.00339f
C6004 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# sky130_fd_sc_hd__conb_1_28/HI -9.78e-19
C6005 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0303f
C6006 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__conb_1_9/LO 7.91e-20
C6007 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.78e-21
C6008 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.303f
C6009 FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_11/Y 7.06e-20
C6010 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_60/Y 2.59e-19
C6011 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_581_47# -7.91e-19
C6012 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.03e-20
C6013 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 1.04e-19
C6014 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_41/HI 9.54e-19
C6015 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 5.83e-19
C6016 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_16_2/Y 0.00986f
C6017 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__conb_1_17/HI 0.0173f
C6018 sky130_fd_sc_hd__conb_1_40/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 6.27e-20
C6019 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_581_47# -2.6e-20
C6020 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# V_LOW -6.55e-19
C6021 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0024f
C6022 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_22/LO 1.81e-20
C6023 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__conb_1_10/HI 2.29e-19
C6024 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__inv_1_61/Y 0.0329f
C6025 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 2.25e-20
C6026 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 1e-20
C6027 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00129f
C6028 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# V_GND -0.00441f
C6029 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_51/Y 0.0368f
C6030 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# V_GND -0.00465f
C6031 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# -9.32e-20
C6032 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_49/LO 4.88e-21
C6033 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# sky130_fd_sc_hd__conb_1_16/HI 2.82e-19
C6034 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# V_LOW 0.0186f
C6035 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 3.22e-19
C6036 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__conb_1_17/HI 2.48e-19
C6037 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__conb_1_12/HI 8.63e-19
C6038 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# -0.00263f
C6039 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# -1.46e-20
C6040 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_557_413# 3.83e-19
C6041 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__conb_1_40/HI 0.0013f
C6042 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 7.93e-21
C6043 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_14/Y 5.78e-20
C6044 sky130_fd_sc_hd__inv_1_98/Y V_LOW 0.101f
C6045 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.37e-19
C6046 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_11/HI 3.23e-20
C6047 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# V_GND -0.00122f
C6048 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__inv_1_103/Y 4.33e-20
C6049 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.578f
C6050 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00161f
C6051 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 5.6e-21
C6052 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# sky130_fd_sc_hd__conb_1_39/HI 2.47e-19
C6053 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 3.04e-19
C6054 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 7.94e-23
C6055 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 0.0044f
C6056 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.35e-20
C6057 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.85e-19
C6058 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.43e-21
C6059 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_103/Y 0.0497f
C6060 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# sky130_fd_sc_hd__conb_1_18/HI 6.25e-20
C6061 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# V_GND 0.00754f
C6062 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# V_GND 0.00625f
C6063 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# -4.66e-20
C6064 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# -3.79e-20
C6065 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# V_LOW 0.0434f
C6066 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 6.3e-19
C6067 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.25e-20
C6068 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 2.11e-19
C6069 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00121f
C6070 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# sky130_fd_sc_hd__conb_1_35/HI 2.05e-19
C6071 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_60/Y 0.211f
C6072 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 3.56e-20
C6073 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 9.14e-19
C6074 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_57/Y 3.07e-20
C6075 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_26/HI 7.81e-20
C6076 Reset sky130_fd_sc_hd__inv_1_63/Y 0.234f
C6077 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 9.4e-21
C6078 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# -0.0285f
C6079 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_557_413# -0.0012f
C6080 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# Reset 1.59e-20
C6081 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__inv_1_47/Y 3.95e-21
C6082 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 4.2e-19
C6083 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00366f
C6084 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0145f
C6085 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 4.32e-20
C6086 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__conb_1_27/LO 3.14e-20
C6087 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.54e-19
C6088 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_85/Y 0.0132f
C6089 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_23/Y 1.89e-19
C6090 sky130_fd_sc_hd__inv_1_95/A Reset 5.37e-19
C6091 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_1_58/Y 3.82e-19
C6092 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# -6.43e-20
C6093 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# -3.06e-20
C6094 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__conb_1_35/HI 0.00741f
C6095 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00164f
C6096 sky130_fd_sc_hd__nand3_1_1/a_109_47# Reset 4.63e-20
C6097 sky130_fd_sc_hd__dfbbn_1_2/Q_N V_GND -0.00686f
C6098 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0163f
C6099 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 3.28e-20
C6100 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# sky130_fd_sc_hd__conb_1_38/HI -6.57e-19
C6101 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__conb_1_29/LO 5.43e-20
C6102 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# V_GND 0.00228f
C6103 sky130_fd_sc_hd__conb_1_36/HI V_GND -0.144f
C6104 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__conb_1_12/LO 1.47e-19
C6105 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_55/Y 0.00503f
C6106 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 7.67e-19
C6107 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/Q_N -4.78e-20
C6108 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# 1.22e-22
C6109 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_63/Y 0.0014f
C6110 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__conb_1_34/LO 3.82e-21
C6111 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 6.36e-19
C6112 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# -3.79e-20
C6113 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# -4.66e-20
C6114 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__conb_1_17/HI 0.0024f
C6115 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 2.66e-20
C6116 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_86/Y 1.03e-19
C6117 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.44e-21
C6118 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 2.48e-19
C6119 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__conb_1_48/HI 0.118f
C6120 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/Q_N -4.16e-20
C6121 RISING_COUNTER.COUNT_SUB_DFF1.Q V_GND 2.09f
C6122 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# sky130_fd_sc_hd__inv_1_55/Y 5.11e-19
C6123 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# -0.00108f
C6124 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__conb_1_46/LO 9.95e-20
C6125 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.36e-20
C6126 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_21/Y 0.0454f
C6127 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# V_LOW -0.00121f
C6128 sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# V_LOW 2.94e-20
C6129 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_16_2/Y 1.12e-19
C6130 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0.00193f
C6131 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# -9.32e-20
C6132 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 3.7e-19
C6133 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__conb_1_12/HI -1.84e-19
C6134 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__inv_1_57/Y 0.00227f
C6135 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__conb_1_40/HI 1.76e-19
C6136 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.0378f
C6137 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 7.48e-19
C6138 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 8.02e-21
C6139 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 7.48e-19
C6140 sky130_fd_sc_hd__inv_1_64/A RISING_COUNTER.COUNT_SUB_DFF5.Q 8.57e-20
C6141 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.14e-20
C6142 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# sky130_fd_sc_hd__inv_1_103/Y 2.07e-20
C6143 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_16_1/Y 0.0538f
C6144 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_44/A 0.147f
C6145 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__inv_1_18/Y 0.00501f
C6146 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 7.44e-19
C6147 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 9.13e-20
C6148 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# Reset 0.00382f
C6149 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.13e-21
C6150 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 1.98e-21
C6151 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF12.Q 1.31e-20
C6152 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0185f
C6153 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# V_GND 0.0209f
C6154 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_54/Y 0.0218f
C6155 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/Q_N -4.78e-20
C6156 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_58/Y 0.192f
C6157 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_557_413# 0.00219f
C6158 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF15.Q 5.69e-19
C6159 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# V_GND 0.00172f
C6160 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0235f
C6161 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# V_GND 7.34e-19
C6162 sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# V_LOW 2.94e-20
C6163 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_71/Y 1.3e-19
C6164 sky130_fd_sc_hd__dfbbn_1_22/a_1363_47# sky130_fd_sc_hd__conb_1_32/HI -6.57e-19
C6165 sky130_fd_sc_hd__conb_1_10/HI V_GND -0.121f
C6166 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_941_21# 0.303f
C6167 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 4.76e-21
C6168 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 2.1e-20
C6169 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.13f
C6170 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_107/Y 0.25f
C6171 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__nand3_1_2/Y 2.47e-20
C6172 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_37/LO 1.04e-20
C6173 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.83e-20
C6174 sky130_fd_sc_hd__inv_1_104/Y V_LOW 0.0129f
C6175 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_1_4/a_113_47# 2.11e-21
C6176 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 5.27e-19
C6177 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__conb_1_7/HI 1.19e-20
C6178 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__conb_1_0/HI 0.00682f
C6179 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# V_GND 0.0079f
C6180 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_103/Y 0.133f
C6181 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_19/HI 0.00195f
C6182 RISING_COUNTER.COUNT_SUB_DFF5.Q V_GND 1.35f
C6183 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 1.02e-21
C6184 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_35/HI 0.0436f
C6185 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# Reset 0.0188f
C6186 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# Reset 6.96e-19
C6187 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# 3.12e-21
C6188 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_1_61/Y 0.00182f
C6189 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_61/Y 2.42e-19
C6190 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# V_GND -0.00153f
C6191 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# CLOCK_GEN.SR_Op.Q 7.03e-21
C6192 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__conb_1_34/HI 0.0198f
C6193 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.48e-19
C6194 sky130_fd_sc_hd__conb_1_5/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 4.53e-21
C6195 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.61e-20
C6196 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00133f
C6197 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0293f
C6198 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.42e-21
C6199 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__conb_1_11/HI 1.16e-20
C6200 sky130_fd_sc_hd__nand2_1_3/Y V_GND -0.00276f
C6201 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_39/HI 0.0615f
C6202 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0341f
C6203 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__inv_1_12/Y 8.88e-19
C6204 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -3.85e-19
C6205 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_891_329# -0.0016f
C6206 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_97/A 3.24e-20
C6207 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.24e-21
C6208 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00164f
C6209 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 6.4e-20
C6210 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.44e-19
C6211 sky130_fd_sc_hd__inv_1_32/Y V_SENSE 0.102f
C6212 sky130_fd_sc_hd__conb_1_10/LO V_LOW 0.102f
C6213 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.0245f
C6214 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_581_47# -2.6e-20
C6215 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 1.13e-19
C6216 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# V_LOW -0.00121f
C6217 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0252f
C6218 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 0.0012f
C6219 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 3.07e-20
C6220 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/Q_N -4.24e-20
C6221 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__inv_1_57/Y 6.95e-21
C6222 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 0.0416f
C6223 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 2.35e-21
C6224 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 1.51e-20
C6225 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 1.51e-20
C6226 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 2.35e-21
C6227 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_9/LO 4.61e-19
C6228 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__conb_1_40/LO 8.84e-20
C6229 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# sky130_fd_sc_hd__conb_1_5/HI 0.00194f
C6230 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__inv_1_102/Y 0.0503f
C6231 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.00536f
C6232 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 0.0011f
C6233 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 0.0344f
C6234 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# V_LOW -0.0587f
C6235 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_1_5/Y 0.016f
C6236 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_56/Y 0.271f
C6237 sky130_fd_sc_hd__inv_1_71/Y CLOCK_GEN.SR_Op.Q 3.31e-20
C6238 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# V_LOW 4.8e-20
C6239 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_557_413# 5.11e-19
C6240 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 7.32e-19
C6241 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# sky130_fd_sc_hd__conb_1_4/HI 5.03e-19
C6242 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 6.33e-20
C6243 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 0.00122f
C6244 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# V_GND 0.0036f
C6245 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__conb_1_40/LO 1.24e-19
C6246 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# 4.2e-20
C6247 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0391f
C6248 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_58/Y 7.93e-20
C6249 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# 0.00195f
C6250 sky130_fd_sc_hd__conb_1_47/HI V_LOW 0.0676f
C6251 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_105/Y 0.00278f
C6252 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00239f
C6253 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.413f
C6254 sky130_fd_sc_hd__conb_1_19/LO V_GND -0.00527f
C6255 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0011f
C6256 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 0.00184f
C6257 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 7e-20
C6258 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# V_GND -0.00518f
C6259 Reset sky130_fd_sc_hd__conb_1_35/HI 0.113f
C6260 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__conb_1_31/HI 2.87e-19
C6261 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_68/A 5.58e-19
C6262 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__conb_1_1/HI -0.00581f
C6263 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 1.85e-20
C6264 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# 6.91e-20
C6265 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# V_GND -9.19e-19
C6266 sky130_fd_sc_hd__inv_1_22/Y V_LOW 0.156f
C6267 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# sky130_fd_sc_hd__conb_1_36/HI 5.79e-19
C6268 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00123f
C6269 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0056f
C6270 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.76e-20
C6271 sky130_fd_sc_hd__inv_1_76/A V_GND 2.35f
C6272 sky130_fd_sc_hd__conb_1_0/LO V_LOW 0.0956f
C6273 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_11/HI -0.00227f
C6274 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__conb_1_51/HI 4.08e-22
C6275 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_95/A 7.55e-21
C6276 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__inv_1_102/Y 0.0492f
C6277 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 1.46f
C6278 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# sky130_fd_sc_hd__conb_1_34/HI 3.98e-19
C6279 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.89e-19
C6280 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_70/A 0.0185f
C6281 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__conb_1_45/HI 7.93e-21
C6282 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 0.0059f
C6283 FALLING_COUNTER.COUNT_SUB_DFF12.Q V_GND 1.1f
C6284 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__conb_1_51/HI 5.66e-19
C6285 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# Reset 7.9e-20
C6286 sky130_fd_sc_hd__conb_1_47/LO sky130_fd_sc_hd__conb_1_47/HI 7.46e-19
C6287 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.97e-19
C6288 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# -0.00385f
C6289 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.62e-21
C6290 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 2.96e-21
C6291 sky130_fd_sc_hd__nand2_8_9/a_27_47# CLOCK_GEN.SR_Op.Q 0.0453f
C6292 sky130_fd_sc_hd__inv_1_6/Y V_LOW 0.17f
C6293 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# sky130_fd_sc_hd__conb_1_2/HI 2.12e-19
C6294 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_891_329# -0.00159f
C6295 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# -0.00953f
C6296 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00157f
C6297 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_106/Y 1.62e-20
C6298 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 7.41e-19
C6299 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 4.18e-19
C6300 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 1.65e-19
C6301 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 4.56e-21
C6302 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__conb_1_11/HI 2.09e-19
C6303 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_75/A 6.97e-20
C6304 sky130_fd_sc_hd__nand2_1_0/Y V_LOW 0.0503f
C6305 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00242f
C6306 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_1_105/Y 7.52e-20
C6307 sky130_fd_sc_hd__inv_1_13/Y V_GND 0.00586f
C6308 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 0.251f
C6309 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_557_413# 3.09e-21
C6310 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__inv_16_0/Y 0.00682f
C6311 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 4.86e-20
C6312 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 3.31e-22
C6313 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 7.6e-19
C6314 sky130_fd_sc_hd__inv_1_43/Y V_LOW 0.1f
C6315 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__inv_16_0/Y 0.00213f
C6316 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.81e-20
C6317 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00707f
C6318 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_29/Q_N 7.56e-19
C6319 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00325f
C6320 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0162f
C6321 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__inv_1_60/Y 8.87e-19
C6322 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_30/HI 3.76e-19
C6323 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.06e-19
C6324 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.2e-20
C6325 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_381_47# 3.76e-21
C6326 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.31e-20
C6327 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.01e-19
C6328 sky130_fd_sc_hd__dfbbn_1_19/a_1159_47# sky130_fd_sc_hd__conb_1_5/HI 0.00199f
C6329 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.16e-20
C6330 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_15/LO 0.00209f
C6331 sky130_fd_sc_hd__dfbbn_1_30/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.72e-19
C6332 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# 0.0118f
C6333 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 1.11e-21
C6334 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 1.11e-21
C6335 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_24/LO 2.32e-20
C6336 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# V_LOW -9.94e-19
C6337 sky130_fd_sc_hd__inv_1_112/Y V_GND 0.379f
C6338 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 2.51e-21
C6339 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 3.42e-21
C6340 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 2.18e-19
C6341 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 0.00163f
C6342 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 1.44e-20
C6343 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__conb_1_42/HI 1.22e-20
C6344 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_10/LO 8.84e-20
C6345 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.12f
C6346 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_647_21# -0.00631f
C6347 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_473_413# -0.00988f
C6348 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_2_0/Y 1.97e-22
C6349 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__inv_1_22/Y 9.63e-19
C6350 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q -4.98e-20
C6351 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__inv_1_99/Y 1.9e-20
C6352 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00517f
C6353 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# V_LOW 0.012f
C6354 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__conb_1_27/HI 8.86e-19
C6355 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0414f
C6356 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_891_329# 8.46e-21
C6357 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 2.96e-19
C6358 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 5.29e-19
C6359 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# V_LOW 0.0288f
C6360 sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__nand3_1_2/Y 3.68e-21
C6361 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.85e-19
C6362 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# 2.47e-21
C6363 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_41/HI 0.0694f
C6364 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# V_LOW 5.38e-19
C6365 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__conb_1_31/HI 2.39e-19
C6366 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# V_GND -3.82e-19
C6367 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_891_329# -2.2e-20
C6368 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_45/HI 0.081f
C6369 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# -0.00751f
C6370 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__conb_1_9/HI -1.02e-19
C6371 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__conb_1_1/HI -1.8e-19
C6372 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__conb_1_36/HI 1.22e-20
C6373 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__inv_1_71/A 2.67e-20
C6374 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 0.00329f
C6375 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0299f
C6376 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__inv_1_22/Y 5.9e-19
C6377 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 1.01e-19
C6378 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_381_47# 3.83e-19
C6379 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 2.03e-21
C6380 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 0.00643f
C6381 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__conb_1_11/HI -2.07e-19
C6382 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0479f
C6383 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_93/Y 0.0024f
C6384 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# V_LOW 0.00493f
C6385 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# V_GND 0.003f
C6386 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_27/LO 8.84e-20
C6387 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# -3.06e-20
C6388 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_647_21# -6.43e-20
C6389 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# V_LOW 8.44e-19
C6390 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# V_GND 0.00875f
C6391 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# V_LOW 0.0295f
C6392 sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# sky130_fd_sc_hd__conb_1_45/HI 4.22e-19
C6393 sky130_fd_sc_hd__dfbbn_1_44/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 2.87e-19
C6394 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# V_GND -0.00253f
C6395 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.0725f
C6396 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 5.11e-20
C6397 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__inv_1_10/Y 8.17e-19
C6398 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# V_GND 3.73e-19
C6399 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__conb_1_13/HI -6.61e-19
C6400 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.42e-19
C6401 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_76/A 0.0303f
C6402 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_193_47# -0.0592f
C6403 sky130_fd_sc_hd__inv_1_101/Y sky130_fd_sc_hd__inv_16_1/Y 2.45e-19
C6404 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__inv_1_103/Y 0.0368f
C6405 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_37/HI 4.74e-21
C6406 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/Q_N -6.48e-19
C6407 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# -0.00592f
C6408 sky130_fd_sc_hd__dfbbn_1_19/Q_N FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00389f
C6409 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.32e-19
C6410 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 2.91e-19
C6411 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 5.13e-19
C6412 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 0.00303f
C6413 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0.00244f
C6414 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 4.39e-20
C6415 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 3.13e-19
C6416 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 0.0312f
C6417 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# Reset 0.00223f
C6418 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__inv_1_108/Y 4.58e-20
C6419 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.19f
C6420 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.19e-20
C6421 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# V_GND 5.27e-19
C6422 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# V_GND 0.00699f
C6423 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# V_LOW 0.0565f
C6424 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 2.12e-19
C6425 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# V_GND 3.31e-19
C6426 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_1_112/Y 0.0235f
C6427 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__inv_1_21/Y 0.00164f
C6428 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# V_LOW -0.0159f
C6429 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.24e-19
C6430 sky130_fd_sc_hd__inv_1_60/Y sky130_fd_sc_hd__conb_1_28/HI 2.37e-19
C6431 transmission_gate_0/GN V_SENSE 0.0313f
C6432 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 0.00286f
C6433 sky130_fd_sc_hd__conb_1_13/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 2.16e-20
C6434 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# V_LOW -0.00602f
C6435 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# V_GND 0.00552f
C6436 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.07e-19
C6437 FALLING_COUNTER.COUNT_SUB_DFF4.Q V_GND 0.6f
C6438 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 3.74e-19
C6439 sky130_fd_sc_hd__conb_1_18/LO V_GND -0.0053f
C6440 sky130_fd_sc_hd__conb_1_37/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0624f
C6441 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.72e-20
C6442 sky130_fd_sc_hd__conb_1_44/HI V_LOW 0.202f
C6443 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_101/Y 0.0626f
C6444 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# -3.48e-20
C6445 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_891_329# -2.2e-20
C6446 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 7.4e-19
C6447 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# Reset 0.0343f
C6448 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__inv_1_62/Y 4.78e-20
C6449 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 4.18e-20
C6450 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 9.07e-21
C6451 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 5.9e-20
C6452 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 2.93e-20
C6453 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 6.21e-20
C6454 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/Q_N 0.0365f
C6455 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 7.62e-20
C6456 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/Q_N 7.62e-20
C6457 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 0.0175f
C6458 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# V_GND -8.43e-19
C6459 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0.598f
C6460 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# sky130_fd_sc_hd__conb_1_22/HI 1.06e-20
C6461 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# V_GND 0.00678f
C6462 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0192f
C6463 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# 9.79e-21
C6464 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 2.82e-20
C6465 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__conb_1_42/HI -6.57e-19
C6466 RISING_COUNTER.COUNT_SUB_DFF4.Q V_LOW 4.28f
C6467 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# -8.61e-20
C6468 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# V_GND 0.00429f
C6469 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_27/LO 1.02e-20
C6470 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0477f
C6471 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# V_GND 2.54e-19
C6472 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__conb_1_20/HI 0.159f
C6473 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0779f
C6474 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# V_LOW 1.79e-20
C6475 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# V_LOW 2.26e-20
C6476 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.466f
C6477 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__conb_1_27/HI 0.00262f
C6478 sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__inv_1_78/A 0.00438f
C6479 sky130_fd_sc_hd__nand2_8_3/Y sky130_fd_sc_hd__inv_1_76/A 0.226f
C6480 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# V_LOW -6.55e-19
C6481 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# -0.0078f
C6482 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# -0.0152f
C6483 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_1_75/A 9.42e-21
C6484 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__inv_1_12/Y 0.132f
C6485 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# V_LOW 2.42e-19
C6486 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__conb_1_31/HI 4.34e-20
C6487 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.0086f
C6488 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.0086f
C6489 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 4.4e-20
C6490 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 4.4e-20
C6491 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_1_20/Y 1.55e-20
C6492 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# -3.46e-20
C6493 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 1.42e-32
C6494 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__conb_1_1/HI -2.17e-19
C6495 sky130_fd_sc_hd__dfbbn_1_46/a_1363_47# sky130_fd_sc_hd__conb_1_36/HI -4.57e-19
C6496 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__conb_1_48/LO 8.84e-20
C6497 sky130_fd_sc_hd__inv_1_79/A V_GND 0.0619f
C6498 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# V_LOW -0.00326f
C6499 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# V_LOW 0.018f
C6500 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__conb_1_47/HI 0.00487f
C6501 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_16_1/Y 0.00124f
C6502 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__inv_1_22/Y 0.0109f
C6503 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 0.00321f
C6504 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# V_GND 0.00432f
C6505 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.81e-19
C6506 sky130_fd_sc_hd__inv_1_65/Y V_LOW 0.151f
C6507 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_1_12/Y 6.15e-19
C6508 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__inv_1_64/A 0.00168f
C6509 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__conb_1_13/HI 1.51e-21
C6510 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_47/Y 0.00583f
C6511 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# V_LOW -1.39e-35
C6512 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# V_GND 1.72e-19
C6513 sky130_fd_sc_hd__nand3_1_2/a_109_47# V_LOW -6.68e-21
C6514 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__inv_1_12/Y 0.00101f
C6515 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# V_GND 0.00194f
C6516 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# V_LOW 0.00836f
C6517 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.7e-20
C6518 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# -0.00813f
C6519 sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# V_GND 5.79e-19
C6520 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.9e-19
C6521 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 4.01e-19
C6522 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 3.03e-19
C6523 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 6.71e-20
C6524 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 5.87e-21
C6525 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 0.00173f
C6526 sky130_fd_sc_hd__conb_1_29/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 1.74e-19
C6527 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__inv_1_9/Y 2.93e-20
C6528 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_21/HI 4.13e-20
C6529 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__conb_1_13/HI -2.07e-19
C6530 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# V_LOW 4.8e-20
C6531 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_30/HI 3.85e-20
C6532 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_71/Y 8.9e-19
C6533 sky130_fd_sc_hd__dfbbn_1_32/Q_N Reset 2.78e-19
C6534 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -2.6e-19
C6535 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# -2.02e-19
C6536 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# -5.54e-21
C6537 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 1.46e-19
C6538 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_55/Y 2.71e-20
C6539 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# V_GND 3.13e-19
C6540 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0303f
C6541 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_22/HI 3e-20
C6542 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 1.7e-19
C6543 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__conb_1_11/HI 0.276f
C6544 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# V_GND -0.0439f
C6545 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__conb_1_34/HI 0.00609f
C6546 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 2.67e-20
C6547 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 5.72e-21
C6548 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_71/A 5.74e-21
C6549 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.29e-20
C6550 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_33/HI 0.0115f
C6551 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 1.25e-20
C6552 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 7.97e-20
C6553 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.93e-21
C6554 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# V_LOW 4.8e-20
C6555 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# V_GND 0.0045f
C6556 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.00347f
C6557 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# V_LOW 2.94e-20
C6558 sky130_fd_sc_hd__conb_1_51/LO FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00415f
C6559 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__inv_1_112/Y 0.0708f
C6560 sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# V_LOW -6.55e-19
C6561 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.82e-19
C6562 sky130_fd_sc_hd__inv_1_88/Y V_GND 0.0434f
C6563 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.03e-21
C6564 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# V_GND -0.151f
C6565 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.86e-20
C6566 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# 5.17e-20
C6567 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# V_LOW 1.04e-19
C6568 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.9e-19
C6569 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# V_GND 2.58e-19
C6570 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# Reset 2.48e-20
C6571 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 6.25e-20
C6572 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# V_GND 0.00232f
C6573 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__conb_1_41/HI 0.00557f
C6574 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0283f
C6575 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_46/LO 2.63e-20
C6576 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 1.04e-20
C6577 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# -3.46e-20
C6578 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.0313f
C6579 sky130_fd_sc_hd__conb_1_51/LO V_LOW 0.0439f
C6580 sky130_fd_sc_hd__dfbbn_1_38/Q_N FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00578f
C6581 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_557_413# -3.67e-20
C6582 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_891_329# -2.46e-19
C6583 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# -0.0279f
C6584 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_18/HI 3.58e-20
C6585 sky130_fd_sc_hd__dfbbn_1_29/a_581_47# Reset 6.07e-19
C6586 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 1.61e-20
C6587 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 2.81e-20
C6588 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# V_GND 1.73e-19
C6589 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0411f
C6590 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.203f
C6591 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# sky130_fd_sc_hd__inv_1_21/Y 1.12e-20
C6592 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# V_GND 6.59e-19
C6593 sky130_fd_sc_hd__inv_1_8/Y V_LOW 0.259f
C6594 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_50/A 0.067f
C6595 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_581_47# -7.91e-19
C6596 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# V_GND 7.25e-19
C6597 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0197f
C6598 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# -0.00149f
C6599 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_101/Y 1.57e-21
C6600 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# V_LOW -0.00266f
C6601 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 7.44e-19
C6602 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 9.13e-20
C6603 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_1_19/Y 6.31e-21
C6604 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# -0.00364f
C6605 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 9.78e-19
C6606 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0.00738f
C6607 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 1.03e-19
C6608 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 1.03e-19
C6609 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 9.78e-19
C6610 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00205f
C6611 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_6/HI 0.00256f
C6612 sky130_fd_sc_hd__nor2_1_0/Y V_LOW 0.21f
C6613 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00641f
C6614 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_39/HI 0.00913f
C6615 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 1.17e-21
C6616 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_83/Y 6.9e-21
C6617 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_473_413# -3.06e-20
C6618 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_647_21# -0.00631f
C6619 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.122f
C6620 sky130_fd_sc_hd__dfbbn_1_34/Q_N V_LOW -0.00396f
C6621 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 3.29e-19
C6622 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 3.29e-19
C6623 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 3.69e-20
C6624 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_791_47# 3.69e-20
C6625 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.00299f
C6626 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.00299f
C6627 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0.00378f
C6628 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_18/Y 0.0336f
C6629 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 8.46e-19
C6630 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__inv_1_102/Y 0.00185f
C6631 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# V_LOW -2.78e-35
C6632 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# 3.53e-19
C6633 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# V_GND -8.97e-19
C6634 FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_16_1/Y 0.207f
C6635 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.55e-19
C6636 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 5.16e-20
C6637 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 7.71e-21
C6638 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__conb_1_13/HI 6.08e-21
C6639 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 5.47e-21
C6640 sky130_fd_sc_hd__dfbbn_1_29/Q_N V_LOW -0.00501f
C6641 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# sky130_fd_sc_hd__inv_1_12/Y 0.00105f
C6642 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__inv_1_49/Y -0.00317f
C6643 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.34e-20
C6644 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 4.68e-21
C6645 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.58e-19
C6646 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_891_329# 0.00135f
C6647 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# V_LOW 0.00217f
C6648 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.00228f
C6649 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# -0.00107f
C6650 sky130_fd_sc_hd__dfbbn_1_46/a_557_413# V_LOW 3.56e-20
C6651 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_891_329# 0.00174f
C6652 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.46e-22
C6653 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__conb_1_41/HI -6.91e-20
C6654 sky130_fd_sc_hd__inv_1_102/Y sky130_fd_sc_hd__conb_1_41/HI 2.59e-19
C6655 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__inv_1_72/A 0.00343f
C6656 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.73e-20
C6657 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# -9.32e-20
C6658 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_70/Y 1.12e-19
C6659 sky130_fd_sc_hd__dfbbn_1_23/a_891_329# sky130_fd_sc_hd__conb_1_32/HI 9.76e-19
C6660 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0892f
C6661 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_1_52/Y 9.13e-21
C6662 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 5e-20
C6663 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_40/LO 7.49e-19
C6664 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# V_LOW -0.00266f
C6665 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_34/A 9e-20
C6666 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_1/Y 0.128f
C6667 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# V_GND 3.39e-19
C6668 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00146f
C6669 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_2_0/Y 0.015f
C6670 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__conb_1_34/HI 5.05e-19
C6671 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 0.00175f
C6672 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# 1.63e-19
C6673 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 1.66e-19
C6674 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 3.52e-20
C6675 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__conb_1_41/HI 3.95e-21
C6676 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# -4.66e-20
C6677 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -2.84e-32
C6678 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_381_47# -3.05e-20
C6679 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 6.32e-19
C6680 sky130_fd_sc_hd__dfbbn_1_11/Q_N V_GND -0.00255f
C6681 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# -2.07e-19
C6682 sky130_fd_sc_hd__inv_1_60/Y V_GND 0.048f
C6683 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_19/Y 0.00382f
C6684 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 5.41e-22
C6685 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.77e-19
C6686 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# V_GND 0.00742f
C6687 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# V_LOW 0.0112f
C6688 sky130_fd_sc_hd__conb_1_31/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00126f
C6689 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# V_GND 1.81e-19
C6690 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF12.Q 8.58e-21
C6691 sky130_fd_sc_hd__dfbbn_1_36/Q_N V_LOW -0.00939f
C6692 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_28/HI 2.24e-19
C6693 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.95e-21
C6694 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 5.86e-19
C6695 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.22e-20
C6696 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 2.86e-21
C6697 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 0.00132f
C6698 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 0.00202f
C6699 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.00221f
C6700 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00103f
C6701 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# V_GND -8.76e-19
C6702 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# sky130_fd_sc_hd__conb_1_41/HI 2.78e-21
C6703 sky130_fd_sc_hd__inv_1_44/A V_GND 0.0803f
C6704 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_17/HI 5.41e-20
C6705 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__conb_1_50/LO 7.48e-20
C6706 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# 4.53e-19
C6707 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -0.00133f
C6708 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# -3.04e-19
C6709 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.00169f
C6710 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 5.05e-19
C6711 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 0.00122f
C6712 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.00106f
C6713 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 4.66e-19
C6714 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_97/A 0.164f
C6715 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# -4.66e-20
C6716 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# V_GND 0.00268f
C6717 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_51/HI 0.00141f
C6718 sky130_fd_sc_hd__inv_1_58/Y V_LOW 0.00675f
C6719 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00109f
C6720 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_581_47# -2.6e-20
C6721 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# 1.07e-19
C6722 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__inv_1_76/A 9.92e-21
C6723 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 0.0011f
C6724 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# V_LOW 0.0241f
C6725 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 0.0143f
C6726 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_1_12/Y 1.24e-21
C6727 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0.00272f
C6728 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# sky130_fd_sc_hd__inv_1_19/Y 9.44e-20
C6729 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_581_47# -2.6e-20
C6730 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 4.01e-20
C6731 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 4.01e-20
C6732 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_16/HI 4.6e-20
C6733 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 3.68e-20
C6734 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 6.78e-19
C6735 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 1.33e-20
C6736 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 1.11e-19
C6737 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 4.54e-19
C6738 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 2.27f
C6739 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0549f
C6740 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# V_LOW -0.108f
C6741 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0427f
C6742 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_21/HI 0.0783f
C6743 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# -0.00344f
C6744 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# -1.61e-19
C6745 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_13/LO 3.6e-19
C6746 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# sky130_fd_sc_hd__inv_1_102/Y 1.57e-19
C6747 sky130_fd_sc_hd__nand2_8_4/a_27_47# Reset 0.0213f
C6748 sky130_fd_sc_hd__dfbbn_1_1/Q_N V_LOW -0.0104f
C6749 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# V_LOW 0.0127f
C6750 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__inv_1_13/Y 2.24e-19
C6751 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__conb_1_36/HI 6.45e-19
C6752 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__inv_1_8/Y 0.00469f
C6753 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_71/A 0.0221f
C6754 sky130_fd_sc_hd__inv_16_2/Y V_GND 3.27f
C6755 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 8.28e-20
C6756 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# V_GND 0.00511f
C6757 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# V_LOW 0.00563f
C6758 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00167f
C6759 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00497f
C6760 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_35/LO 0.00841f
C6761 sky130_fd_sc_hd__inv_1_70/Y CLOCK_GEN.SR_Op.Q 4.59e-20
C6762 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 1.2e-21
C6763 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 0.0156f
C6764 sky130_fd_sc_hd__inv_1_101/Y V_LOW 0.168f
C6765 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 6.21e-21
C6766 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.08e-20
C6767 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.45e-19
C6768 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__inv_1_53/Y 2.28e-19
C6769 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# V_GND -0.0051f
C6770 sky130_fd_sc_hd__conb_1_1/HI Reset 7.38e-19
C6771 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 2.65e-19
C6772 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 0.00236f
C6773 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/Q_N -4.24e-20
C6774 sky130_fd_sc_hd__fill_4_73/VPB V_LOW 0.797f
C6775 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# V_GND 0.00539f
C6776 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_70/Y 8.86e-20
C6777 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# V_GND 0.00631f
C6778 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 7.63e-19
C6779 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 7.63e-19
C6780 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_18/LO 5.7e-21
C6781 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# sky130_fd_sc_hd__inv_1_15/Y 4.63e-20
C6782 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.29e-19
C6783 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_46/a_381_47# 2.04e-21
C6784 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 6.29e-19
C6785 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_27_47# -0.00307f
C6786 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 9.94e-20
C6787 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__inv_1_103/Y 2.39e-19
C6788 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# V_GND -0.00858f
C6789 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_1_108/Y 3.97e-19
C6790 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# -0.00336f
C6791 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_16/Y 0.00139f
C6792 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_381_47# -3.79e-20
C6793 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_1_12/Y 0.23f
C6794 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# V_LOW 2.94e-20
C6795 sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__inv_1_61/Y 0.025f
C6796 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.92e-20
C6797 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_16_0/Y 2.84e-19
C6798 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__inv_1_7/Y 0.00111f
C6799 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.59e-21
C6800 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 0.00519f
C6801 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 7.01e-21
C6802 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 1.28f
C6803 sky130_fd_sc_hd__dfbbn_1_32/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00164f
C6804 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_35/HI 0.00301f
C6805 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 5.01e-19
C6806 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 0.00707f
C6807 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 2.23e-21
C6808 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 8.17e-21
C6809 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 3.84e-21
C6810 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0241f
C6811 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 0.0133f
C6812 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.395f
C6813 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 4.17e-20
C6814 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 5.29e-19
C6815 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0167f
C6816 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_1_23/Y -2.87e-20
C6817 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00141f
C6818 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_35/a_381_47# 4.4e-19
C6819 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 6.05e-20
C6820 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.425f
C6821 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# V_GND -0.00155f
C6822 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_50/A 0.00214f
C6823 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_43/A 2.05e-21
C6824 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__conb_1_51/HI 6.95e-21
C6825 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 4.6e-20
C6826 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 4.64e-20
C6827 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 3.79e-19
C6828 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 5.67e-20
C6829 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0.00401f
C6830 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0.00334f
C6831 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 3.22e-19
C6832 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 9.08e-19
C6833 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 3.88e-19
C6834 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# V_LOW 2.94e-20
C6835 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 2.62e-20
C6836 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.03e-19
C6837 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# 3.72e-19
C6838 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__conb_1_33/LO 3.14e-20
C6839 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.0062f
C6840 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 5.45e-19
C6841 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# 1.08e-20
C6842 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__conb_1_23/HI 1.72e-20
C6843 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_110/Y 1.97e-20
C6844 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0901f
C6845 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0302f
C6846 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 9.71e-20
C6847 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0.00117f
C6848 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 9.56e-19
C6849 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 1.67e-20
C6850 RISING_COUNTER.COUNT_SUB_DFF7.Q V_LOW 1.66f
C6851 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__conb_1_46/HI -0.00119f
C6852 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# V_LOW -8.84e-19
C6853 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__conb_1_2/HI 0.028f
C6854 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0294f
C6855 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0025f
C6856 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# -2.57e-20
C6857 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__conb_1_13/LO 9.83e-21
C6858 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__inv_1_103/Y 0.00109f
C6859 sky130_fd_sc_hd__inv_1_104/Y FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.008f
C6860 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_59/Y 0.00749f
C6861 Reset sky130_fd_sc_hd__inv_1_90/Y 0.0169f
C6862 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 3.47e-21
C6863 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_35/LO 1.68e-19
C6864 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# V_LOW 1.51e-20
C6865 sky130_fd_sc_hd__nand2_1_2/a_113_47# V_LOW -1.78e-19
C6866 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_100/Y 2.74e-19
C6867 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_15/Y 0.00906f
C6868 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 9.69e-21
C6869 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# V_GND 7.25e-19
C6870 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.00372f
C6871 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.24e-19
C6872 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0274f
C6873 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1_23/HI 0.00206f
C6874 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# 0.0048f
C6875 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.00218f
C6876 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 9.69e-20
C6877 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 1.3e-19
C6878 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 4.45e-20
C6879 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_64/A 5.12e-19
C6880 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.0018f
C6881 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 0.00349f
C6882 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__inv_1_102/Y 1.56e-21
C6883 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_26/LO 8.84e-20
C6884 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 1.25e-19
C6885 FALLING_COUNTER.COUNT_SUB_DFF3.Q V_GND 0.628f
C6886 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# V_LOW 0.0176f
C6887 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 2.02e-22
C6888 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 3.95e-21
C6889 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 2.39e-20
C6890 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 2.16e-20
C6891 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 3.6e-21
C6892 sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# V_GND -3.7e-19
C6893 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_20/Y 7.8e-20
C6894 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00359f
C6895 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 4.43e-20
C6896 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 0.00106f
C6897 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.013f
C6898 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00466f
C6899 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0287f
C6900 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.0029f
C6901 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# V_GND 2.72e-19
C6902 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.33e-20
C6903 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# -6.22e-19
C6904 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# -0.00538f
C6905 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# -6.23e-21
C6906 sky130_fd_sc_hd__fill_4_84/VPB V_GND 0.393f
C6907 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# V_GND 0.00399f
C6908 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_941_21# 0.00175f
C6909 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 2.76e-19
C6910 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# 2.76e-19
C6911 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_97/Y 0.0215f
C6912 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 0.0016f
C6913 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 0.00514f
C6914 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 0.0016f
C6915 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 0.00514f
C6916 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 3.58e-20
C6917 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.422f
C6918 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# V_GND -0.185f
C6919 sky130_fd_sc_hd__conb_1_19/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 2.14e-19
C6920 sky130_fd_sc_hd__conb_1_5/LO sky130_fd_sc_hd__conb_1_5/HI 0.00126f
C6921 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# V_GND -0.0203f
C6922 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# -3.79e-20
C6923 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# -0.00336f
C6924 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -9.31e-20
C6925 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.26f
C6926 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 9.6e-21
C6927 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__inv_1_47/Y 1.31e-20
C6928 sky130_fd_sc_hd__inv_1_96/A V_GND 0.215f
C6929 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# V_GND 0.009f
C6930 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__conb_1_35/HI 5.45e-20
C6931 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 3.15e-19
C6932 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# sky130_fd_sc_hd__conb_1_45/HI 5.72e-19
C6933 sky130_fd_sc_hd__conb_1_29/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0916f
C6934 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.19e-21
C6935 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 1.83e-21
C6936 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/Q_N -9.56e-20
C6937 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.21e-20
C6938 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.94e-19
C6939 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.35e-20
C6940 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.00101f
C6941 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_791_47# 1.4e-20
C6942 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_108/Y 0.00483f
C6943 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.82e-19
C6944 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.25e-21
C6945 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# V_GND 0.0152f
C6946 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0363f
C6947 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_92/Y 1.04e-20
C6948 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_647_21# 2.83e-20
C6949 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00616f
C6950 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_91/A 4.43e-21
C6951 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00526f
C6952 CLOCK_GEN.SR_Op.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 2.19f
C6953 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_16_0/Y 2.65e-19
C6954 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.87e-20
C6955 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.14f
C6956 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 5.85e-19
C6957 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_1_18/Y 7.05e-20
C6958 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 6.57e-19
C6959 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.27e-20
C6960 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.0187f
C6961 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 4.13e-20
C6962 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_23/Y 1.71e-21
C6963 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0436f
C6964 sky130_fd_sc_hd__dfbbn_1_8/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 9.23e-19
C6965 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 5.38e-19
C6966 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 6.28e-21
C6967 sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 7.49e-20
C6968 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# sky130_fd_sc_hd__conb_1_24/HI 4.78e-20
C6969 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__conb_1_33/HI 0.00398f
C6970 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# sky130_fd_sc_hd__conb_1_46/HI 8.63e-19
C6971 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# sky130_fd_sc_hd__conb_1_2/HI 2.22e-20
C6972 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# -8.96e-20
C6973 sky130_fd_sc_hd__dfbbn_1_33/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00209f
C6974 FALLING_COUNTER.COUNT_SUB_DFF9.Q V_LOW 1.04f
C6975 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# -4.37e-20
C6976 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# -6.23e-21
C6977 sky130_fd_sc_hd__conb_1_7/LO V_LOW 0.0966f
C6978 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_12/HI 0.137f
C6979 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI 0.00517f
C6980 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_1_20/Y 0.00506f
C6981 sky130_fd_sc_hd__inv_1_55/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 5.78e-20
C6982 sky130_fd_sc_hd__conb_1_25/LO V_GND -0.00511f
C6983 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_71/A 5.04e-20
C6984 sky130_fd_sc_hd__conb_1_32/LO V_GND 0.00155f
C6985 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.00364f
C6986 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# V_GND -0.155f
C6987 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.287f
C6988 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 8.98e-21
C6989 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 3.79e-20
C6990 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/Q_N 0.00814f
C6991 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 0.00294f
C6992 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 0.00156f
C6993 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 2.26e-20
C6994 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# sky130_fd_sc_hd__conb_1_45/HI 3.53e-19
C6995 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# V_LOW 3.56e-20
C6996 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# V_LOW -0.00174f
C6997 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.06e-21
C6998 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_76/A 1.96e-19
C6999 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 3.11e-19
C7000 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# V_LOW 0.00609f
C7001 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__inv_1_99/Y 5.91e-20
C7002 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 1.13e-20
C7003 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# -2.74e-21
C7004 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# -0.00263f
C7005 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__inv_1_100/Y 4.54e-19
C7006 sky130_fd_sc_hd__conb_1_43/LO V_GND -0.00405f
C7007 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00226f
C7008 sky130_fd_sc_hd__dfbbn_1_39/a_557_413# sky130_fd_sc_hd__inv_16_1/Y 0.00214f
C7009 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# V_LOW -9.15e-19
C7010 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_0/HI 4.84e-20
C7011 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_16/HI 0.0377f
C7012 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__inv_1_22/Y 0.0134f
C7013 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# 1.04e-19
C7014 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 2.02e-19
C7015 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.13e-19
C7016 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.87e-20
C7017 sky130_fd_sc_hd__conb_1_47/LO FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.08e-19
C7018 sky130_fd_sc_hd__dfbbn_1_3/Q_N V_GND 4.12e-19
C7019 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00482f
C7020 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 3.01e-20
C7021 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_791_47# 3.01e-20
C7022 sky130_fd_sc_hd__dfbbn_1_18/a_557_413# V_LOW 3.56e-20
C7023 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 9.87e-21
C7024 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# V_GND 1.42e-19
C7025 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# V_GND 2.54e-19
C7026 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# sky130_fd_sc_hd__conb_1_22/HI 8.54e-20
C7027 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# V_LOW 0.0329f
C7028 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_557_413# -3.67e-20
C7029 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# -5.33e-20
C7030 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_891_329# 0.00285f
C7031 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# V_GND 1.44e-19
C7032 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_2/LO 5.26e-19
C7033 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# V_GND 3.46e-19
C7034 sky130_fd_sc_hd__inv_1_31/A V_GND 0.0214f
C7035 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_17/HI 1.36e-20
C7036 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# V_GND 1.12e-19
C7037 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# V_LOW 0.016f
C7038 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF9.Q 7.9e-19
C7039 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_5/LO 0.00422f
C7040 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -0.0115f
C7041 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# -2.28e-19
C7042 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_11/HI 0.00916f
C7043 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 1.84e-19
C7044 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.0141f
C7045 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 3.24e-21
C7046 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_70/Y 2.43e-19
C7047 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00284f
C7048 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__conb_1_26/HI 1.46e-19
C7049 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# -2.37e-19
C7050 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -0.0116f
C7051 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# 6.83e-21
C7052 sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# V_GND 1.39e-19
C7053 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__conb_1_22/HI 0.0377f
C7054 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0589f
C7055 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__inv_1_59/Y 9.75e-19
C7056 sky130_fd_sc_hd__dfbbn_1_44/a_557_413# V_GND 2.59e-19
C7057 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0322f
C7058 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 3.65e-20
C7059 sky130_fd_sc_hd__conb_1_3/HI V_LOW 0.139f
C7060 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0426f
C7061 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__conb_1_42/HI 8.97e-21
C7062 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# Reset 2.47e-19
C7063 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00119f
C7064 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0144f
C7065 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.16f
C7066 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_95/A 5.96e-20
C7067 sky130_fd_sc_hd__inv_1_9/Y V_GND 0.031f
C7068 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 0.0158f
C7069 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.52e-19
C7070 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_21/a_27_47# 0.0118f
C7071 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__inv_1_18/Y 4.7e-20
C7072 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# V_LOW 3.56e-20
C7073 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# V_GND 0.00489f
C7074 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 2.09e-20
C7075 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# -0.00548f
C7076 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 4.15e-19
C7077 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00106f
C7078 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_41/HI 5.21e-20
C7079 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_1_65/Y 0.0238f
C7080 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 3.92e-22
C7081 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 3.92e-22
C7082 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_94/A 0.0147f
C7083 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00359f
C7084 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# sky130_fd_sc_hd__conb_1_33/HI -5.73e-20
C7085 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.79e-20
C7086 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -5.54e-21
C7087 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -2.18e-19
C7088 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1_70/Y 0.00507f
C7089 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# sky130_fd_sc_hd__inv_1_21/Y 2.81e-19
C7090 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 8.86e-21
C7091 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 3.31e-19
C7092 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.92e-19
C7093 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_90/Y 0.00112f
C7094 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# -0.00548f
C7095 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_891_329# -0.00159f
C7096 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__inv_1_60/Y 3.42e-20
C7097 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# V_GND 8.77e-20
C7098 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# V_LOW -2.78e-35
C7099 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# sky130_fd_sc_hd__inv_1_17/Y 0.00156f
C7100 sky130_fd_sc_hd__nand3_1_2/B V_GND 0.313f
C7101 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0275f
C7102 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__conb_1_8/HI 3.11e-20
C7103 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 3.1e-20
C7104 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__conb_1_38/LO 1.33e-19
C7105 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# -9.32e-20
C7106 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# sky130_fd_sc_hd__inv_1_100/Y 2.34e-19
C7107 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0474f
C7108 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# V_LOW -3.49e-19
C7109 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__conb_1_50/LO 1.53e-19
C7110 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_17/HI 3.28e-20
C7111 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 7.14e-19
C7112 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 8.51e-19
C7113 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_25/HI 0.0233f
C7114 sky130_fd_sc_hd__conb_1_33/LO sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 8.84e-20
C7115 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_83/Y 1.8e-19
C7116 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0413f
C7117 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 9.4e-20
C7118 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# V_LOW 0.016f
C7119 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# sky130_fd_sc_hd__inv_1_105/Y 7.09e-19
C7120 sky130_fd_sc_hd__inv_2_0/A transmission_gate_0/GN 0.00119f
C7121 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.99e-20
C7122 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# V_GND 0.0126f
C7123 sky130_fd_sc_hd__inv_1_102/Y V_GND 0.189f
C7124 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.501f
C7125 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# -0.00149f
C7126 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.92e-19
C7127 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# V_GND 3.04e-19
C7128 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# -1.64e-19
C7129 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_12/LO 5e-20
C7130 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.108f
C7131 FULL_COUNTER.COUNT_SUB_DFF13.Q V_GND 1.15f
C7132 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0.00378f
C7133 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.81e-20
C7134 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 9.03e-19
C7135 sky130_fd_sc_hd__inv_1_49/Y V_GND 0.111f
C7136 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1e-18
C7137 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# sky130_fd_sc_hd__conb_1_26/HI 8.79e-21
C7138 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# -0.00985f
C7139 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_647_21# -0.00631f
C7140 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# -7.17e-20
C7141 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# -1.66e-19
C7142 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 0.0144f
C7143 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_72/A 1.43e-20
C7144 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 7.41e-19
C7145 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.89e-20
C7146 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_2/Y 0.02f
C7147 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_3/Y 0.0112f
C7148 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.935f
C7149 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0559f
C7150 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 3.12e-19
C7151 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_35/LO 4.53e-21
C7152 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# sky130_fd_sc_hd__conb_1_42/HI 1.29e-20
C7153 sky130_fd_sc_hd__dfbbn_1_31/a_581_47# Reset 6.71e-20
C7154 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00334f
C7155 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.79e-19
C7156 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 2.48e-19
C7157 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 5.71e-19
C7158 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# V_GND 0.0105f
C7159 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_21/a_27_47# 2.33e-19
C7160 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00216f
C7161 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_891_329# -0.00159f
C7162 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# -0.014f
C7163 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__conb_1_38/HI 4.95e-19
C7164 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# V_GND 2.56e-19
C7165 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__inv_16_0/Y 0.434f
C7166 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_581_47# -2.6e-20
C7167 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_16_0/Y 0.0044f
C7168 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__conb_1_41/HI 1.07e-20
C7169 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__conb_1_20/HI 0.00419f
C7170 FULL_COUNTER.COUNT_SUB_DFF8.Q V_LOW 1.01f
C7171 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 4.57e-19
C7172 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.37e-20
C7173 sky130_fd_sc_hd__conb_1_33/LO Reset 0.00403f
C7174 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__conb_1_33/HI -2.17e-19
C7175 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 0.00132f
C7176 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0.00132f
C7177 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 3.9e-19
C7178 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.34e-22
C7179 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_12/Y 4.85e-21
C7180 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_20/Y 1.27e-19
C7181 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 8.91e-20
C7182 sky130_fd_sc_hd__inv_1_78/A sky130_fd_sc_hd__inv_1_97/Y 0.0376f
C7183 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# -1.03e-19
C7184 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# -3.86e-20
C7185 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 6.55e-19
C7186 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_941_21# 0.0211f
C7187 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_4/LO 6.57e-20
C7188 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# -0.00171f
C7189 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF3.Q 4.87e-20
C7190 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# -3.46e-20
C7191 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00101f
C7192 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00314f
C7193 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 4.13e-19
C7194 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# -0.0166f
C7195 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_891_329# -2.2e-20
C7196 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 5.08e-19
C7197 sky130_fd_sc_hd__dfbbn_1_26/Q_N V_LOW -0.00509f
C7198 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_46/A 0.0346f
C7199 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.92e-20
C7200 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__conb_1_8/HI 7.51e-20
C7201 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_647_21# 9.61e-19
C7202 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.68e-19
C7203 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# V_LOW -0.00266f
C7204 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_891_329# -0.00161f
C7205 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# -0.00524f
C7206 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.93e-19
C7207 sky130_fd_sc_hd__dfbbn_1_31/Q_N V_LOW -0.0011f
C7208 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.00359f
C7209 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/Q_N -4.24e-20
C7210 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 2.45e-19
C7211 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 1.42e-19
C7212 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 6.61e-19
C7213 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__conb_1_24/HI 0.00173f
C7214 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_68/A 0.0253f
C7215 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.38e-21
C7216 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_76/A 0.032f
C7217 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 7.5e-19
C7218 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 7.5e-20
C7219 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.77e-21
C7220 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.63e-21
C7221 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.46e-22
C7222 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 6.08e-21
C7223 sky130_fd_sc_hd__conb_1_32/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 1.46e-20
C7224 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_70/A 0.0314f
C7225 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__inv_1_90/Y 0.0107f
C7226 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__conb_1_25/HI 6.18e-20
C7227 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.96e-19
C7228 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__inv_1_9/Y 2.91e-21
C7229 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# V_GND -0.133f
C7230 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 0.17f
C7231 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0434f
C7232 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 9.79e-21
C7233 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_25/LO 0.0103f
C7234 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# V_GND -8.97e-19
C7235 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__inv_1_99/Y 2.57e-19
C7236 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.366f
C7237 sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 0.00286f
C7238 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# V_LOW 4.8e-20
C7239 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 3.3e-20
C7240 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_581_47# -2.6e-20
C7241 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 0.107f
C7242 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 1.96e-19
C7243 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_106/Y 2.68e-20
C7244 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_1_104/Y 4.09e-22
C7245 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0.303f
C7246 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.93e-20
C7247 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00914f
C7248 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 4.53e-19
C7249 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 3.5e-19
C7250 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 6.96e-21
C7251 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.139f
C7252 sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 0.00129f
C7253 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 7.06e-21
C7254 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.09e-19
C7255 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.36e-20
C7256 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# sky130_fd_sc_hd__inv_1_19/Y 0.00103f
C7257 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__inv_1_59/Y 2.22e-20
C7258 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# 1.24e-19
C7259 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0411f
C7260 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 8.69e-19
C7261 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.298f
C7262 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__inv_1_61/Y 5.2e-20
C7263 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 5.53e-21
C7264 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# 2.87e-19
C7265 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# V_GND 2.47e-19
C7266 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_100/Y 0.022f
C7267 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# -0.00592f
C7268 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__conb_1_28/HI 4.15e-21
C7269 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__conb_1_6/HI 6.56e-21
C7270 sky130_fd_sc_hd__dfbbn_1_20/a_581_47# sky130_fd_sc_hd__conb_1_20/HI 6.07e-19
C7271 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00786f
C7272 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 2.86e-19
C7273 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 2.7e-20
C7274 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 7.35e-21
C7275 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.05e-19
C7276 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 8.12e-21
C7277 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 7.74e-19
C7278 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_110/Y 7.29e-20
C7279 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# -2.57e-20
C7280 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/Q_N -4.33e-20
C7281 sky130_fd_sc_hd__inv_1_18/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0195f
C7282 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_11/HI 0.423f
C7283 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 6.52e-22
C7284 sky130_fd_sc_hd__inv_1_74/Y V_GND 0.263f
C7285 sky130_fd_sc_hd__nand3_1_2/B sky130_fd_sc_hd__nand2_8_3/Y 4.6e-19
C7286 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_93/A 2.31e-19
C7287 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.11e-19
C7288 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 7.35e-19
C7289 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 5.79e-19
C7290 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.00182f
C7291 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# -1.44e-20
C7292 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.17e-20
C7293 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/Q_N -6.48e-19
C7294 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_581_47# 5.8e-19
C7295 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.06e-19
C7296 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 2.91e-20
C7297 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# -0.00592f
C7298 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00349f
C7299 CLOCK_GEN.SR_Op.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00226f
C7300 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 2.46e-19
C7301 sky130_fd_sc_hd__dfbbn_1_39/a_557_413# V_LOW -9.15e-19
C7302 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__inv_1_53/Y 0.00259f
C7303 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 8.33e-21
C7304 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.07e-19
C7305 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__conb_1_8/HI 2.05e-19
C7306 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# -0.00385f
C7307 sky130_fd_sc_hd__dfbbn_1_28/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 1.12e-19
C7308 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0449f
C7309 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__conb_1_8/HI 4.04e-19
C7310 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# 4.84e-19
C7311 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_53/Y 0.0396f
C7312 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00264f
C7313 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 4.03e-21
C7314 sky130_fd_sc_hd__dfbbn_1_19/Q_N V_LOW -0.00505f
C7315 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# CLOCK_GEN.SR_Op.Q 5.65e-21
C7316 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00102f
C7317 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__inv_1_8/Y 2.1e-19
C7318 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.3e-19
C7319 sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__conb_1_13/HI 5.94e-20
C7320 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# CLOCK_GEN.SR_Op.Q 0.0297f
C7321 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# V_LOW 3.13e-19
C7322 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 2.91e-21
C7323 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.91e-22
C7324 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 0.00324f
C7325 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0.00493f
C7326 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0628f
C7327 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__conb_1_12/HI 4.28e-21
C7328 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__inv_1_9/Y 1.17e-22
C7329 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# V_GND 1.25e-19
C7330 FULL_COUNTER.COUNT_SUB_DFF0.Q V_LOW 8.04f
C7331 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_105/Y 2.29e-20
C7332 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00137f
C7333 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00691f
C7334 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 9.65e-20
C7335 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_1_11/Y 5.93e-20
C7336 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 9.42e-19
C7337 sky130_fd_sc_hd__inv_1_81/Y V_LOW 0.421f
C7338 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 0.002f
C7339 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.22e-20
C7340 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.4e-19
C7341 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.05e-19
C7342 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.65e-20
C7343 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0397f
C7344 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# 7.17e-19
C7345 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.08e-20
C7346 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 9.18e-19
C7347 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 9.03e-21
C7348 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# V_GND 0.0124f
C7349 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_381_47# 3.76e-19
C7350 FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_6/HI 0.308f
C7351 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_1_112/Y 2.54e-23
C7352 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0589f
C7353 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 3.35e-19
C7354 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__conb_1_42/HI 0.00196f
C7355 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_97/Y 0.104f
C7356 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 0.0174f
C7357 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_21/LO 5.04e-21
C7358 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__conb_1_28/LO 5.27e-20
C7359 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 4.91e-21
C7360 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__conb_1_21/HI 0.00138f
C7361 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_16/HI 0.0933f
C7362 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 4.31e-19
C7363 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 1.16e-19
C7364 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 3.59e-19
C7365 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__nand3_1_1/a_193_47# 5.15e-20
C7366 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 2.11e-21
C7367 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 6.36e-19
C7368 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 0.00284f
C7369 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_473_413# -3.06e-20
C7370 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_647_21# -6.43e-20
C7371 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 6.27e-20
C7372 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_14/LO 0.0093f
C7373 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_0/HI 0.0119f
C7374 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_98/Y 0.382f
C7375 sky130_fd_sc_hd__inv_1_52/Y V_GND 0.195f
C7376 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_44/A 0.00152f
C7377 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 4.57e-19
C7378 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__conb_1_34/LO 1.33e-19
C7379 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 3.51e-21
C7380 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 0.0013f
C7381 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.02e-19
C7382 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 0.00116f
C7383 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00126f
C7384 sky130_fd_sc_hd__dfbbn_1_30/Q_N FALLING_COUNTER.COUNT_SUB_DFF1.Q 4.49e-20
C7385 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_72/A 0.0351f
C7386 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# sky130_fd_sc_hd__conb_1_25/HI 5.67e-19
C7387 sky130_fd_sc_hd__dfbbn_1_8/Q_N FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0363f
C7388 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0397f
C7389 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 7.28e-21
C7390 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# sky130_fd_sc_hd__inv_1_101/Y 7.09e-19
C7391 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 0.0253f
C7392 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_26/HI 0.0323f
C7393 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_12/HI 0.0133f
C7394 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__conb_1_30/HI 0.00943f
C7395 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# -4.43e-19
C7396 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# -3.86e-20
C7397 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_45/LO 8.84e-20
C7398 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.36e-21
C7399 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.77e-20
C7400 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 4.98e-20
C7401 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_7/HI 0.0697f
C7402 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_72/A 0.00308f
C7403 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 1.59e-19
C7404 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.98e-19
C7405 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__conb_1_5/LO 0.00168f
C7406 sky130_fd_sc_hd__inv_1_119/Y sky130_fd_sc_hd__inv_1_76/A 0.376f
C7407 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.43e-20
C7408 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.43e-20
C7409 sky130_fd_sc_hd__dfbbn_1_28/a_891_329# sky130_fd_sc_hd__inv_1_54/Y 4.87e-19
C7410 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_1_76/A 0.00155f
C7411 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__conb_1_39/HI 3.89e-21
C7412 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 3.7e-19
C7413 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_38/Q_N 5.2e-20
C7414 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 6.03e-19
C7415 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.78e-19
C7416 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.32e-19
C7417 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 2.47e-20
C7418 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# V_LOW 0.00623f
C7419 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00598f
C7420 sky130_fd_sc_hd__conb_1_6/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 1.95e-19
C7421 sky130_fd_sc_hd__inv_1_59/Y V_GND 0.0846f
C7422 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# 0.00632f
C7423 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 7.48e-21
C7424 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00482f
C7425 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_647_21# -0.00431f
C7426 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# -0.0105f
C7427 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.91e-19
C7428 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# V_GND 0.00453f
C7429 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.66e-19
C7430 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.05f
C7431 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_23/Y 3.74e-20
C7432 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00147f
C7433 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 0.00507f
C7434 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_50/Y 2.01e-19
C7435 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0215f
C7436 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 1.51e-19
C7437 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# CLOCK_GEN.SR_Op.Q 2.66e-20
C7438 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.16e-19
C7439 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# V_LOW 0.0185f
C7440 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# V_GND 0.00438f
C7441 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.335f
C7442 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0026f
C7443 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# V_GND 0.0106f
C7444 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# V_LOW 0.0205f
C7445 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 9.87e-19
C7446 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__nand2_8_3/Y 1.59e-19
C7447 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_94/A 4.05e-24
C7448 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__conb_1_19/LO 0.0551f
C7449 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 4.94e-19
C7450 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# V_GND 0.00318f
C7451 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.37e-19
C7452 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# V_LOW 0.0146f
C7453 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_37/LO 2.38e-19
C7454 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.66e-20
C7455 sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# sky130_fd_sc_hd__conb_1_21/HI 1.79e-19
C7456 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF8.Q 0.372f
C7457 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.09e-21
C7458 sky130_fd_sc_hd__inv_1_1/Y V_SENSE 0.466f
C7459 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 2.66e-19
C7460 sky130_fd_sc_hd__dfbbn_1_35/Q_N sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 8.22e-20
C7461 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_891_329# -0.00159f
C7462 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# -0.00947f
C7463 sky130_fd_sc_hd__conb_1_45/LO sky130_fd_sc_hd__conb_1_44/HI 8.84e-20
C7464 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_30/HI 1.93e-20
C7465 sky130_fd_sc_hd__conb_1_34/LO RISING_COUNTER.COUNT_SUB_DFF4.Q 1.16e-19
C7466 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.37e-21
C7467 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_1_6/Y 1.07e-20
C7468 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_1_107/Y 8.75e-21
C7469 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0279f
C7470 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 4e-20
C7471 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00146f
C7472 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__inv_1_98/Y 0.00641f
C7473 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_16_1/Y 1.24e-20
C7474 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# V_GND 0.00434f
C7475 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# V_GND 0.00433f
C7476 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.45e-19
C7477 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 0.0012f
C7478 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 0.00413f
C7479 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# V_GND 0.00651f
C7480 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 7.93e-21
C7481 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 1.07e-20
C7482 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00791f
C7483 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_891_329# 0.00119f
C7484 sky130_fd_sc_hd__conb_1_27/LO RISING_COUNTER.COUNT_SUB_DFF2.Q 0.139f
C7485 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__conb_1_28/HI 0.00209f
C7486 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_44/HI 0.00592f
C7487 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__nand3_1_0/Y 0.0415f
C7488 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__conb_1_16/HI 1.34e-19
C7489 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__inv_1_106/Y 0.00127f
C7490 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# -6.23e-21
C7491 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# -0.00367f
C7492 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# -0.00631f
C7493 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# -0.00985f
C7494 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__conb_1_16/HI 0.00115f
C7495 sky130_fd_sc_hd__dfbbn_1_26/a_581_47# sky130_fd_sc_hd__conb_1_30/HI 1.52e-19
C7496 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# -2.57e-20
C7497 sky130_fd_sc_hd__nand3_1_0/Y V_GND 0.0962f
C7498 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 1.3e-19
C7499 sky130_fd_sc_hd__dfbbn_1_43/Q_N RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00668f
C7500 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_647_21# -0.00122f
C7501 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# -0.00312f
C7502 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__conb_1_51/HI 3.12e-19
C7503 sky130_fd_sc_hd__dfbbn_1_6/a_1363_47# sky130_fd_sc_hd__conb_1_10/HI -4.57e-19
C7504 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# V_LOW -0.315f
C7505 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_557_413# 0.00156f
C7506 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 3.31e-21
C7507 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 1.02e-21
C7508 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.07e-19
C7509 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# V_GND -7.73e-19
C7510 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__conb_1_18/HI 1.16e-20
C7511 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__inv_16_1/Y 0.429f
C7512 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# sky130_fd_sc_hd__conb_1_22/HI 3.32e-19
C7513 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# V_GND -8.97e-19
C7514 sky130_fd_sc_hd__inv_1_51/A V_GND 0.147f
C7515 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# -9.88e-20
C7516 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# -0.00175f
C7517 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# -0.00199f
C7518 sky130_fd_sc_hd__inv_1_94/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 1.01e-24
C7519 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_1_18/Y 2.47e-20
C7520 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 3.07e-20
C7521 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.91e-20
C7522 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.0106f
C7523 sky130_fd_sc_hd__conb_1_17/HI V_LOW 0.106f
C7524 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.29e-20
C7525 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__conb_1_48/HI 5.47e-20
C7526 sky130_fd_sc_hd__dfbbn_1_42/a_557_413# V_LOW 3.56e-20
C7527 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__conb_1_12/HI 7.93e-21
C7528 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# 0.00808f
C7529 sky130_fd_sc_hd__nand2_8_2/A V_GND 0.141f
C7530 sky130_fd_sc_hd__conb_1_16/HI FULL_COUNTER.COUNT_SUB_DFF18.Q 1.68e-19
C7531 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_47/Y 0.0623f
C7532 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# V_LOW -0.00266f
C7533 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 8.08e-21
C7534 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_32/HI 0.0717f
C7535 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 4.06e-21
C7536 sky130_fd_sc_hd__dfbbn_1_21/Q_N V_GND 0.00369f
C7537 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# V_GND -0.0453f
C7538 sky130_fd_sc_hd__conb_1_37/HI Reset 0.0311f
C7539 FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_11/Y 2.87e-20
C7540 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.04e-19
C7541 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__conb_1_39/HI 0.00487f
C7542 sky130_fd_sc_hd__dfbbn_1_50/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 5.48e-19
C7543 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# CLOCK_GEN.SR_Op.Q 2.23e-19
C7544 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# 5.39e-19
C7545 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.62e-19
C7546 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# CLOCK_GEN.SR_Op.Q 9.94e-21
C7547 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_1_18/Y 0.0548f
C7548 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# -3.04e-19
C7549 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# -6.23e-21
C7550 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 6.66e-19
C7551 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# V_LOW 1.79e-20
C7552 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__inv_1_57/Y 0.00226f
C7553 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# 9.1e-21
C7554 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# V_GND 0.00143f
C7555 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00177f
C7556 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# -0.208f
C7557 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00503f
C7558 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF1.Q 4.39e-19
C7559 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# V_GND 1.58e-19
C7560 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00233f
C7561 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_35/HI 0.00514f
C7562 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# V_GND -9.03e-19
C7563 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_54/Y 5.81e-20
C7564 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__conb_1_40/HI 9.82e-19
C7565 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_32/LO 0.00221f
C7566 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 5.23e-19
C7567 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 9.16e-20
C7568 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 5.37e-19
C7569 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 1.01e-19
C7570 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__conb_1_40/HI 0.00306f
C7571 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.07e-20
C7572 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.3e-19
C7573 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00625f
C7574 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0329f
C7575 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__conb_1_9/HI 1.32e-20
C7576 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# -0.00592f
C7577 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0119f
C7578 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.42e-20
C7579 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0546f
C7580 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI 1.23e-19
C7581 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.03e-20
C7582 FALLING_COUNTER.COUNT_SUB_DFF10.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 1f
C7583 sky130_fd_sc_hd__inv_1_75/Y V_LOW 0.285f
C7584 sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# V_GND 3.24e-19
C7585 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 1e-19
C7586 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 3.74e-20
C7587 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 2.37e-20
C7588 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# V_GND -0.00211f
C7589 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__nand3_1_2/B 0.0459f
C7590 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# V_LOW 4.8e-20
C7591 Reset sky130_fd_sc_hd__inv_1_93/A 0.0457f
C7592 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nand3_1_1/Y 0.184f
C7593 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 0.00613f
C7594 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# V_GND 0.00519f
C7595 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 2.3e-20
C7596 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# V_LOW -0.00266f
C7597 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_941_21# 6.94e-19
C7598 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_16_1/Y 0.395f
C7599 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_45/HI 3.65e-19
C7600 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_9/LO 4.39e-19
C7601 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.43e-21
C7602 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0559f
C7603 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.81e-20
C7604 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 3.12e-19
C7605 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_193_47# -0.23f
C7606 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__conb_1_17/HI 0.00244f
C7607 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__conb_1_40/HI 4.9e-19
C7608 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00119f
C7609 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 1.68e-21
C7610 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# V_GND -9.27e-19
C7611 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.44e-20
C7612 sky130_fd_sc_hd__dfbbn_1_7/Q_N FULL_COUNTER.COUNT_SUB_DFF17.Q 5.25e-19
C7613 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00222f
C7614 sky130_fd_sc_hd__dfbbn_1_47/a_581_47# V_GND -9.08e-19
C7615 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_100/Y 0.362f
C7616 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__inv_16_0/Y 0.0101f
C7617 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0223f
C7618 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# 3.42e-20
C7619 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 0.0105f
C7620 sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 2.66e-19
C7621 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 4.69e-21
C7622 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# V_LOW 0.0226f
C7623 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_8/HI 2.07e-20
C7624 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# -0.00827f
C7625 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# -0.00125f
C7626 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__conb_1_17/HI 2.13e-19
C7627 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# sky130_fd_sc_hd__conb_1_12/HI -4.09e-19
C7628 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_891_329# 0.00144f
C7629 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# sky130_fd_sc_hd__conb_1_40/HI 5.21e-19
C7630 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/Q_N 0.0015f
C7631 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_11/HI 6.87e-19
C7632 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 0.213f
C7633 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# V_GND 2.36e-19
C7634 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0314f
C7635 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__conb_1_16/HI 4.12e-20
C7636 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.177f
C7637 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_47/HI 0.0574f
C7638 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# sky130_fd_sc_hd__conb_1_39/HI -0.00185f
C7639 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.13e-20
C7640 RISING_COUNTER.COUNT_SUB_DFF0.Q V_LOW 1.18f
C7641 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0.00372f
C7642 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_1_17/Y 3.55e-19
C7643 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# sky130_fd_sc_hd__inv_1_18/Y 0.00101f
C7644 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.21e-19
C7645 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 6.89e-21
C7646 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# 6.95e-21
C7647 sky130_fd_sc_hd__dfbbn_1_37/Q_N V_GND 0.00151f
C7648 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# V_GND 0.005f
C7649 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# V_GND 0.00152f
C7650 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.37e-19
C7651 sky130_fd_sc_hd__dfbbn_1_13/Q_N FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0306f
C7652 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# V_LOW 0.0106f
C7653 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 4.39e-20
C7654 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.003f
C7655 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.37e-20
C7656 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_112/Y 0.0718f
C7657 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 3.74e-20
C7658 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# -0.00796f
C7659 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_891_329# -0.00159f
C7660 FALLING_COUNTER.COUNT_SUB_DFF5.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00465f
C7661 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 3.64e-19
C7662 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 4.32e-21
C7663 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 4.07e-19
C7664 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.043f
C7665 sky130_fd_sc_hd__conb_1_23/LO RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00216f
C7666 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_10/LO 0.00126f
C7667 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 3.58e-20
C7668 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__conb_1_27/LO 2.6e-19
C7669 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_1_6/Y 5.85e-22
C7670 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00359f
C7671 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_72/A 0.0013f
C7672 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -9.35e-20
C7673 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# -3.86e-20
C7674 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_58/Y 1.07e-21
C7675 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 1.05e-20
C7676 sky130_fd_sc_hd__nand3_1_1/a_193_47# Reset 2.12e-19
C7677 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__conb_1_35/HI 1.96e-19
C7678 sky130_fd_sc_hd__nand2_8_3/a_27_47# V_LOW -0.00931f
C7679 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# V_GND -0.0464f
C7680 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__conb_1_29/LO 2.76e-21
C7681 sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__conb_1_30/HI 2.07e-20
C7682 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0.013f
C7683 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_67/Y 4.54e-19
C7684 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0411f
C7685 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# 3.62e-21
C7686 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 0.00224f
C7687 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__inv_1_63/Y 1.1e-20
C7688 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 0.00137f
C7689 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# CLOCK_GEN.SR_Op.Q 5.46e-19
C7690 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00328f
C7691 sky130_fd_sc_hd__dfbbn_1_12/a_581_47# sky130_fd_sc_hd__conb_1_17/HI 0.00211f
C7692 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 5.98e-19
C7693 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/Q_N 3.32e-20
C7694 sky130_fd_sc_hd__conb_1_23/HI V_GND -0.228f
C7695 sky130_fd_sc_hd__nand2_8_3/Y sky130_fd_sc_hd__nand2_8_2/A 0.00839f
C7696 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_67/Y 1.77e-19
C7697 sky130_fd_sc_hd__conb_1_25/HI V_GND -0.0365f
C7698 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00118f
C7699 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__conb_1_48/HI 0.041f
C7700 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/Q_N -9.56e-20
C7701 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# sky130_fd_sc_hd__inv_1_55/Y 5.11e-19
C7702 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 8.04e-19
C7703 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 3.56e-19
C7704 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# -3.06e-20
C7705 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# -0.00631f
C7706 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.49e-20
C7707 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# V_LOW -0.00266f
C7708 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 3.45e-20
C7709 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_1_57/Y 0.0017f
C7710 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 0.0199f
C7711 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 2.85e-19
C7712 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 2.85e-19
C7713 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0027f
C7714 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 3.88e-19
C7715 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 5.94e-19
C7716 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 4.12e-19
C7717 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_26/HI 0.00195f
C7718 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_1_102/Y 1.41e-19
C7719 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# 2.26e-21
C7720 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# V_LOW 0.0267f
C7721 sky130_fd_sc_hd__fill_4_85/VPB V_LOW 0.798f
C7722 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_11/LO 0.059f
C7723 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# sky130_fd_sc_hd__inv_1_100/Y 2.2e-21
C7724 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0397f
C7725 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# V_GND 0.00922f
C7726 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_891_329# 0.00289f
C7727 sky130_fd_sc_hd__inv_1_104/Y FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0161f
C7728 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_98/Y 0.107f
C7729 sky130_fd_sc_hd__dfbbn_1_33/a_581_47# V_GND 2.58e-19
C7730 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 1.02e-19
C7731 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_53/Y 2.04e-19
C7732 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# V_GND 3.11e-19
C7733 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0178f
C7734 sky130_fd_sc_hd__fill_4_72/VPB V_GND 0.392f
C7735 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.3e-22
C7736 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.35e-21
C7737 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# 0.113f
C7738 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 9.42e-21
C7739 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 2.28e-20
C7740 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_107/Y 0.294f
C7741 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# -0.00282f
C7742 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__conb_1_41/HI 0.0116f
C7743 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__nand3_1_2/Y 0.0165f
C7744 sky130_fd_sc_hd__dfbbn_1_26/Q_N RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0326f
C7745 sky130_fd_sc_hd__inv_1_71/A V_LOW 1.46f
C7746 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__conb_1_0/HI 0.0028f
C7747 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand3_1_2/Y 9.99e-19
C7748 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 1.7e-19
C7749 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# V_GND -0.00256f
C7750 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_103/Y 0.166f
C7751 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# -2.57e-20
C7752 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_19/HI 2.28e-20
C7753 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# Reset 0.0118f
C7754 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__conb_1_35/HI 1.69e-19
C7755 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# Reset 1.5e-19
C7756 sky130_fd_sc_hd__dfbbn_1_21/Q_N RISING_COUNTER.COUNT_SUB_DFF12.Q 8.63e-19
C7757 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__inv_1_61/Y 0.00571f
C7758 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_61/Y 2.47e-19
C7759 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# CLOCK_GEN.SR_Op.Q 1.22e-20
C7760 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# V_GND 2.47e-19
C7761 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__conb_1_34/HI 0.00521f
C7762 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.3e-19
C7763 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_57/Y 4.56e-21
C7764 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0297f
C7765 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.85e-21
C7766 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_93/A 1.71e-19
C7767 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__inv_1_59/Y 3.47e-19
C7768 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# CLOCK_GEN.SR_Op.Q 2.82e-20
C7769 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_24/HI 0.00541f
C7770 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.0102f
C7771 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.344f
C7772 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0202f
C7773 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# 9.44e-20
C7774 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_10/a_381_47# -3.79e-20
C7775 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# -0.00336f
C7776 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__conb_1_34/LO 2.18e-20
C7777 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 1.19e-19
C7778 sky130_fd_sc_hd__inv_1_105/Y V_GND 0.236f
C7779 sky130_fd_sc_hd__conb_1_42/HI V_LOW 0.0903f
C7780 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 3.77e-19
C7781 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0.00421f
C7782 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.144f
C7783 sky130_fd_sc_hd__conb_1_3/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 2.62e-19
C7784 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_80/A 1.71e-19
C7785 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.488f
C7786 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 3.83e-20
C7787 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 3.45e-20
C7788 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__conb_1_48/HI 0.0494f
C7789 CLOCK_GEN.SR_Op.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 4.06e-21
C7790 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 0.0704f
C7791 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 2.54e-20
C7792 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__conb_1_41/HI 6.46e-19
C7793 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 3.93e-20
C7794 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# V_LOW -0.00266f
C7795 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0111f
C7796 sky130_fd_sc_hd__conb_1_43/HI RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00133f
C7797 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/Q_N -9.56e-20
C7798 Reset transmission_gate_0/GN 0.0488f
C7799 sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# sky130_fd_sc_hd__inv_16_1/Y 0.00113f
C7800 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF2.Q 9.95e-19
C7801 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__conb_1_9/LO 6.63e-19
C7802 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 0.0038f
C7803 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0088f
C7804 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__inv_1_67/Y 0.00133f
C7805 sky130_fd_sc_hd__dfbbn_1_39/Q_N sky130_fd_sc_hd__inv_1_103/Y 1.6e-20
C7806 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 4.97e-20
C7807 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_791_47# 1.03e-20
C7808 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# V_LOW -0.00709f
C7809 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_381_47# 7.13e-22
C7810 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_22/HI 4.68e-19
C7811 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# V_LOW 2.94e-20
C7812 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_891_329# 5.1e-19
C7813 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__inv_1_98/Y 7.39e-19
C7814 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# sky130_fd_sc_hd__conb_1_4/HI 0.00134f
C7815 sky130_fd_sc_hd__inv_1_102/Y sky130_fd_sc_hd__inv_1_100/Y 1.04e-19
C7816 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_1_13/Y 2.23e-21
C7817 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0635f
C7818 sky130_fd_sc_hd__dfbbn_1_28/a_581_47# V_GND 4.43e-19
C7819 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 6.02e-19
C7820 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 0.0124f
C7821 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.00799f
C7822 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__inv_1_76/A 1.04e-19
C7823 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF7.Q 1.2f
C7824 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 9.87e-21
C7825 sky130_fd_sc_hd__dfbbn_1_27/a_581_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00271f
C7826 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_58/Y 4.32e-20
C7827 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_31/Y 0.0959f
C7828 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_31/A 4.69e-19
C7829 FULL_COUNTER.COUNT_SUB_DFF3.Q V_GND 0.598f
C7830 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# 0.0356f
C7831 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_1_105/Y 0.0112f
C7832 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 1.54e-20
C7833 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# sky130_fd_sc_hd__inv_1_107/Y 0.00885f
C7834 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.0546f
C7835 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00172f
C7836 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__dfbbn_1_37/Q_N 3.01e-19
C7837 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 6.17e-20
C7838 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__conb_1_31/HI 0.0205f
C7839 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# V_GND 1.72e-19
C7840 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_10/HI 0.00331f
C7841 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__inv_16_2/Y 0.103f
C7842 sky130_fd_sc_hd__inv_1_92/Y Reset 0.0285f
C7843 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# sky130_fd_sc_hd__conb_1_0/HI 1.79e-19
C7844 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__conb_1_1/HI 1.22e-20
C7845 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_76/A 0.125f
C7846 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# V_GND -0.00164f
C7847 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__inv_1_103/Y 0.00386f
C7848 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# sky130_fd_sc_hd__conb_1_36/HI 0.00211f
C7849 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__conb_1_35/HI 0.00165f
C7850 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# Reset 0.00826f
C7851 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.0406f
C7852 FALLING_COUNTER.COUNT_SUB_DFF6.Q V_LOW 1.12f
C7853 sky130_fd_sc_hd__nand2_1_4/a_113_47# V_LOW -1.78e-19
C7854 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__nand2_1_0/Y 0.215f
C7855 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__conb_1_51/HI 2.06e-19
C7856 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 1.19e-20
C7857 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_11/HI -0.0084f
C7858 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_14/HI 6.77e-19
C7859 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# CLOCK_GEN.SR_Op.Q 4.06e-21
C7860 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# sky130_fd_sc_hd__conb_1_34/HI -1.33e-19
C7861 sky130_fd_sc_hd__inv_1_48/Y FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.285f
C7862 sky130_fd_sc_hd__conb_1_49/LO sky130_fd_sc_hd__conb_1_49/HI 0.00619f
C7863 sky130_fd_sc_hd__fill_4_87/VPB V_LOW 0.797f
C7864 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_67/Y 6.55e-19
C7865 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_40/HI 7.99e-23
C7866 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 3.49e-19
C7867 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 8.65e-20
C7868 sky130_fd_sc_hd__conb_1_26/HI V_LOW 0.0104f
C7869 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_1/Q_N 3.66e-20
C7870 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# -0.00336f
C7871 sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 9.62e-20
C7872 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0.00104f
C7873 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 2.2e-20
C7874 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_85/A 0.222f
C7875 RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0165f
C7876 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_97/A 0.0806f
C7877 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00483f
C7878 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_53/Y 0.24f
C7879 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_1_105/Y 0.0063f
C7880 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__inv_1_53/Y 0.0105f
C7881 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__inv_1_21/Y 0.0361f
C7882 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_891_329# 8.14e-21
C7883 sky130_fd_sc_hd__conb_1_40/HI sky130_fd_sc_hd__conb_1_41/HI 0.0449f
C7884 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 1.47e-20
C7885 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_22/HI 0.0158f
C7886 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_6/HI 0.00527f
C7887 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 1.95e-20
C7888 sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00111f
C7889 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.00269f
C7890 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 1.73e-19
C7891 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__inv_1_57/Y 4.28e-21
C7892 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.87e-19
C7893 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 3.21e-20
C7894 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/Q_N 3.21e-20
C7895 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.11e-20
C7896 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.23e-19
C7897 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_24/LO 2.57e-19
C7898 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# 4.63e-19
C7899 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# V_LOW 0.00147f
C7900 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_22/HI 3.18e-20
C7901 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 4.82e-19
C7902 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.721f
C7903 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0425f
C7904 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_941_21# -0.00215f
C7905 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_473_413# -0.0103f
C7906 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF12.Q 1.08f
C7907 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__inv_1_22/Y 0.00279f
C7908 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.69e-19
C7909 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# V_LOW 0.0188f
C7910 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF12.Q 7e-20
C7911 sky130_fd_sc_hd__inv_1_62/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 2.1e-19
C7912 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_68/A 0.00335f
C7913 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__conb_1_27/HI 0.00249f
C7914 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# sky130_fd_sc_hd__inv_1_105/Y 0.0255f
C7915 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# 6.88e-19
C7916 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.42e-19
C7917 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 0.0365f
C7918 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 0.00155f
C7919 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_60/Y -0.00396f
C7920 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# V_LOW -0.311f
C7921 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__conb_1_10/HI 0.00138f
C7922 sky130_fd_sc_hd__inv_1_20/Y V_LOW 0.236f
C7923 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0014f
C7924 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# 2.16e-20
C7925 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# V_LOW -0.00389f
C7926 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# sky130_fd_sc_hd__conb_1_31/HI 5.02e-20
C7927 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# sky130_fd_sc_hd__conb_1_9/HI -0.00221f
C7928 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# -4.66e-20
C7929 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_381_47# -3.79e-20
C7930 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# sky130_fd_sc_hd__conb_1_1/HI -4.57e-19
C7931 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_50/A 0.0107f
C7932 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__conb_1_47/HI 0.00494f
C7933 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__inv_1_22/Y 4.94e-20
C7934 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_941_21# 7.89e-19
C7935 sky130_fd_sc_hd__dfbbn_1_33/Q_N Reset 8.36e-21
C7936 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 7.09e-21
C7937 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 0.00153f
C7938 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 5.52e-20
C7939 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__conb_1_11/HI -0.00118f
C7940 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# V_LOW 1.38e-19
C7941 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# V_GND 4.6e-19
C7942 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# V_GND 0.00648f
C7943 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# -1.61e-20
C7944 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_473_413# -3.86e-20
C7945 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# V_LOW -0.11f
C7946 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# V_LOW 0.00702f
C7947 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 8.55e-19
C7948 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# V_GND 0.0054f
C7949 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.00154f
C7950 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# sky130_fd_sc_hd__inv_1_10/Y 7.05e-19
C7951 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# V_GND 5.57e-19
C7952 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__conb_1_13/HI -0.0076f
C7953 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_647_21# -0.00159f
C7954 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.19e-19
C7955 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# V_LOW 0.0431f
C7956 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_37/HI 3.15e-19
C7957 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 4.26e-21
C7958 sky130_fd_sc_hd__inv_1_70/A V_LOW 0.274f
C7959 sky130_fd_sc_hd__conb_1_44/LO sky130_fd_sc_hd__inv_16_1/Y 0.0373f
C7960 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 6.66e-20
C7961 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 2.88e-19
C7962 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 2.33e-19
C7963 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.01e-19
C7964 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 9.78e-19
C7965 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 1.04e-19
C7966 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.31e-20
C7967 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__nand2_8_0/a_27_47# 0.038f
C7968 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 0.0309f
C7969 FULL_COUNTER.COUNT_SUB_DFF5.Q V_GND 1.37f
C7970 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# Reset 8.37e-19
C7971 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 4.62e-20
C7972 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_71/Y 3.64e-19
C7973 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# V_GND 0.0012f
C7974 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_44/HI 0.164f
C7975 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# V_GND 0.00274f
C7976 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# V_LOW 0.0443f
C7977 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# V_LOW 0.0128f
C7978 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# V_GND 5.14e-19
C7979 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# sky130_fd_sc_hd__inv_1_105/Y 0.0227f
C7980 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# sky130_fd_sc_hd__inv_1_112/Y 0.0014f
C7981 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# V_LOW -0.317f
C7982 sky130_fd_sc_hd__conb_1_21/LO RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0352f
C7983 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.62e-19
C7984 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 7.44e-19
C7985 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 8.44e-20
C7986 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00337f
C7987 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# V_LOW -0.00371f
C7988 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.96e-20
C7989 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# V_GND 0.00298f
C7990 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.76e-19
C7991 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 0.00186f
C7992 sky130_fd_sc_hd__conb_1_17/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00443f
C7993 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.45e-19
C7994 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_101/Y 0.00106f
C7995 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_47/LO 3.51e-20
C7996 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_381_47# -3.79e-20
C7997 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# -4.66e-20
C7998 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 0.0715f
C7999 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.42e-20
C8000 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__conb_1_0/HI 1.86e-19
C8001 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# Reset 0.0246f
C8002 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_66/Y 0.419f
C8003 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 0.00384f
C8004 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 4.07e-19
C8005 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 3.53e-20
C8006 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 4.17e-20
C8007 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.00136f
C8008 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# 8.67e-19
C8009 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.14e-20
C8010 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# V_GND 6.21e-19
C8011 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0.0308f
C8012 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# sky130_fd_sc_hd__conb_1_22/HI 6.86e-20
C8013 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# V_GND 0.00742f
C8014 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_102/Y 0.0405f
C8015 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00157f
C8016 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# 2.83e-19
C8017 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.01e-20
C8018 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# -0.00631f
C8019 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# -0.0109f
C8020 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# V_GND -0.0399f
C8021 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_16_1/Y 0.00825f
C8022 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_12/Y 3.53e-19
C8023 sky130_fd_sc_hd__inv_1_71/Y V_GND 1.11f
C8024 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# V_LOW 0.0293f
C8025 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# V_GND 3.91e-19
C8026 sky130_fd_sc_hd__conb_1_14/LO V_GND -0.00425f
C8027 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 7.69e-20
C8028 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# -9.41e-19
C8029 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__inv_1_53/Y 2.65e-19
C8030 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_58/Y 0.333f
C8031 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_49/Y 0.0292f
C8032 sky130_fd_sc_hd__dfbbn_1_42/a_581_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.86e-19
C8033 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# V_LOW 0.00371f
C8034 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.575f
C8035 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.35e-20
C8036 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0503f
C8037 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# V_LOW 4.8e-20
C8038 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# sky130_fd_sc_hd__conb_1_27/HI 2.13e-19
C8039 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_16_0/Y 1.44e-20
C8040 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 4.26e-20
C8041 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# -0.0225f
C8042 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -0.00415f
C8043 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_86/Y 0.00383f
C8044 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_45/A 0.0291f
C8045 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_7/LO 0.00115f
C8046 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_75/A 6.18e-19
C8047 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__inv_1_20/Y 7.45e-20
C8048 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 0.0149f
C8049 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 7.03e-19
C8050 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.0149f
C8051 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 3.52e-19
C8052 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 7.03e-19
C8053 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 3.52e-19
C8054 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# sky130_fd_sc_hd__conb_1_9/HI -2.07e-19
C8055 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 1.87e-19
C8056 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 3.35e-19
C8057 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# V_LOW -0.00383f
C8058 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF14.Q 4.56e-21
C8059 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# V_LOW 0.0144f
C8060 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# sky130_fd_sc_hd__conb_1_47/HI 6.57e-19
C8061 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# 6.85e-20
C8062 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_193_47# -9.51e-19
C8063 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# V_GND -0.00334f
C8064 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_85/Y 0.0787f
C8065 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.8e-19
C8066 sky130_fd_sc_hd__inv_1_112/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 5.27e-21
C8067 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_1_12/Y 1.56e-19
C8068 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__conb_1_13/HI 3.56e-21
C8069 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__conb_1_11/HI -2.17e-19
C8070 sky130_fd_sc_hd__conb_1_16/LO V_LOW 0.095f
C8071 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# V_LOW -9.94e-19
C8072 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__inv_1_12/Y 0.0392f
C8073 sky130_fd_sc_hd__nand3_1_2/a_193_47# V_LOW -4.49e-19
C8074 sky130_fd_sc_hd__dfbbn_1_20/a_581_47# V_GND 2.66e-19
C8075 sky130_fd_sc_hd__conb_1_23/LO V_LOW 0.0757f
C8076 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# -1.06e-19
C8077 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.2e-20
C8078 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_557_413# -0.0012f
C8079 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# -0.00335f
C8080 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# V_GND 2.24e-19
C8081 sky130_fd_sc_hd__nand2_8_1/a_27_47# V_GND 0.0101f
C8082 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 2.02e-21
C8083 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# 6.25e-21
C8084 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 5.96e-23
C8085 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0128f
C8086 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_581_47# 4.99e-19
C8087 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_1_9/Y 4.41e-21
C8088 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_21/HI 1.39e-19
C8089 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__conb_1_13/HI -3.11e-21
C8090 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_581_47# -7.91e-19
C8091 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.67e-19
C8092 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# V_LOW 2.94e-20
C8093 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# -6.22e-19
C8094 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# -0.00117f
C8095 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# -0.00367f
C8096 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__conb_1_37/HI 1.76e-20
C8097 sky130_fd_sc_hd__inv_1_15/Y V_GND 0.232f
C8098 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# V_GND 4.68e-19
C8099 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.19e-19
C8100 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# V_LOW -0.0189f
C8101 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# V_GND -0.00857f
C8102 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF2.Q 0.43f
C8103 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__conb_1_34/HI 4.72e-19
C8104 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 5.77e-21
C8105 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 2.51e-19
C8106 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 1.05e-20
C8107 sky130_fd_sc_hd__nand2_8_9/a_27_47# V_GND 0.0191f
C8108 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_13/HI 1.35e-19
C8109 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 1.3e-20
C8110 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 1.36e-20
C8111 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.79e-20
C8112 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 5.96e-19
C8113 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_193_47# -0.0818f
C8114 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# sky130_fd_sc_hd__inv_1_108/Y 1.38e-19
C8115 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# V_GND 3.24e-19
C8116 sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# V_LOW 2.94e-20
C8117 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_1_112/Y 3.61e-20
C8118 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# 0.00446f
C8119 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# sky130_fd_sc_hd__conb_1_44/HI 9.76e-19
C8120 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# sky130_fd_sc_hd__inv_1_112/Y 0.0103f
C8121 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.18e-19
C8122 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# V_GND 1.6e-19
C8123 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.21e-20
C8124 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0018f
C8125 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0023f
C8126 sky130_fd_sc_hd__fill_4_68/VPB V_GND 0.382f
C8127 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.25e-19
C8128 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# V_GND 6.75e-19
C8129 sky130_fd_sc_hd__conb_1_33/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 0.227f
C8130 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# Reset 3.66e-19
C8131 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 5.73e-21
C8132 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__nand3_1_1/Y 0.191f
C8133 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_76/A 0.0371f
C8134 Reset sky130_fd_sc_hd__inv_1_67/Y 1.83e-20
C8135 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# V_GND -0.00341f
C8136 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__conb_1_41/HI 0.00568f
C8137 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.0314f
C8138 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_891_329# -2.2e-20
C8139 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# -0.017f
C8140 sky130_fd_sc_hd__inv_1_15/Y sky130_fd_sc_hd__inv_1_12/Y 0.0271f
C8141 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.63e-19
C8142 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 3.78e-19
C8143 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 4.33e-19
C8144 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 7.49e-21
C8145 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# V_GND -0.00153f
C8146 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0479f
C8147 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0724f
C8148 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# V_GND 1.24e-19
C8149 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/Q_N 1.01e-19
C8150 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_8_2/A 2.95e-21
C8151 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_193_47# -0.0319f
C8152 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# V_GND 1.18e-19
C8153 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__inv_1_101/Y 0.00102f
C8154 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# V_LOW -6.55e-19
C8155 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# -3.06e-20
C8156 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_647_21# -6.43e-20
C8157 sky130_fd_sc_hd__dfbbn_1_34/Q_N FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0286f
C8158 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 4.12e-19
C8159 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 5.94e-19
C8160 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 3.88e-19
C8161 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__conb_1_12/HI 0.0168f
C8162 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__conb_1_17/HI 0.0465f
C8163 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# -0.00864f
C8164 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# -0.00312f
C8165 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 7.99e-19
C8166 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 7.99e-19
C8167 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.78e-19
C8168 sky130_fd_sc_hd__dfbbn_1_38/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.73e-19
C8169 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 5.29e-19
C8170 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_23/LO 2.49e-21
C8171 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# -9.41e-19
C8172 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# -0.00408f
C8173 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_473_413# -0.0103f
C8174 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__inv_1_75/A 1.44e-21
C8175 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.033f
C8176 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 6.12e-19
C8177 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_78/A 6.39e-20
C8178 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 6.12e-19
C8179 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.00318f
C8180 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 8.26e-19
C8181 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 8.26e-19
C8182 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 1.1e-19
C8183 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__conb_1_44/HI 0.00139f
C8184 FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_4/Y 6.74e-20
C8185 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__inv_1_102/Y 8.09e-19
C8186 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 8.63e-20
C8187 sky130_fd_sc_hd__conb_1_30/LO V_GND 0.00698f
C8188 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__inv_1_22/Y 1.7e-19
C8189 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_791_47# -0.0127f
C8190 sky130_fd_sc_hd__inv_1_2/Y V_GND 0.0429f
C8191 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# V_GND 7.25e-19
C8192 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.48e-19
C8193 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__conb_1_22/HI 2.73e-22
C8194 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.47e-21
C8195 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 4.66e-22
C8196 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 5.66e-20
C8197 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__conb_1_29/LO 0.00202f
C8198 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__inv_1_49/Y 0.0656f
C8199 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# sky130_fd_sc_hd__inv_1_12/Y 0.00142f
C8200 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.42e-20
C8201 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.48e-20
C8202 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__inv_16_2/Y 1.76e-20
C8203 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 1.25e-19
C8204 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# 0.00202f
C8205 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# V_LOW -7.15e-19
C8206 sky130_fd_sc_hd__dfbbn_1_8/Q_N V_LOW -0.00131f
C8207 sky130_fd_sc_hd__conb_1_41/LO V_GND 0.00252f
C8208 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__nand2_8_3/A 0.152f
C8209 sky130_fd_sc_hd__dfbbn_1_46/a_891_329# V_LOW 2.26e-20
C8210 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# 0.00241f
C8211 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00143f
C8212 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__conb_1_13/HI -2.17e-19
C8213 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__conb_1_41/HI -0.00173f
C8214 sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# sky130_fd_sc_hd__conb_1_32/HI 0.0015f
C8215 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__conb_1_40/LO 1.85e-19
C8216 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00608f
C8217 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# V_LOW -1.01e-19
C8218 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# V_GND -0.0113f
C8219 sky130_fd_sc_hd__conb_1_2/HI V_GND 0.143f
C8220 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 2.21e-19
C8221 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 0.00673f
C8222 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 1.31e-20
C8223 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_19/LO 6.57e-20
C8224 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 6.27e-21
C8225 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 1.13e-19
C8226 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 7.82e-20
C8227 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.213f
C8228 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# -2.92e-20
C8229 sky130_fd_sc_hd__conb_1_27/HI V_LOW 0.0277f
C8230 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00194f
C8231 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# V_GND 0.00797f
C8232 sky130_fd_sc_hd__dfbbn_1_29/Q_N sky130_fd_sc_hd__inv_1_112/Y 0.0248f
C8233 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# -0.205f
C8234 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# V_LOW 0.0109f
C8235 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# V_GND -0.00488f
C8236 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 2.57e-20
C8237 sky130_fd_sc_hd__dfbbn_1_44/Q_N RISING_COUNTER.COUNT_SUB_DFF3.Q 8.95e-21
C8238 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 1.05e-19
C8239 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 8.58e-22
C8240 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 6.27e-20
C8241 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 6.28e-20
C8242 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 3.32e-19
C8243 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.0012f
C8244 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 5.48e-19
C8245 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.98e-20
C8246 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# V_GND -0.00114f
C8247 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__conb_1_41/HI 0.0175f
C8248 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00197f
C8249 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/Q_N -7.11e-33
C8250 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 0.00635f
C8251 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_381_47# -0.00375f
C8252 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# -0.00592f
C8253 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# -1.42e-32
C8254 sky130_fd_sc_hd__inv_1_23/Y V_LOW 0.00688f
C8255 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0.00106f
C8256 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 0.0035f
C8257 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.0029f
C8258 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 0.0034f
C8259 sky130_fd_sc_hd__dfbbn_1_24/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 9.3e-19
C8260 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00173f
C8261 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1_16/HI 1.42e-21
C8262 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_1_22/Y 3.64e-19
C8263 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_39/A 1.93e-19
C8264 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# V_GND -0.0447f
C8265 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__conb_1_51/HI 0.00173f
C8266 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_381_47# 0.00348f
C8267 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__inv_1_76/A 7.07e-20
C8268 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 4.97e-20
C8269 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_791_47# 1.03e-20
C8270 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# V_LOW 0.0143f
C8271 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_80/A 0.0319f
C8272 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_557_413# 0.0022f
C8273 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 2.76e-19
C8274 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_1_12/Y 5.93e-19
C8275 sky130_fd_sc_hd__inv_1_88/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.08f
C8276 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0124f
C8277 sky130_fd_sc_hd__inv_1_103/Y V_GND 0.233f
C8278 sky130_fd_sc_hd__inv_1_19/Y sky130_fd_sc_hd__conb_1_11/HI 0.0528f
C8279 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 3.01e-20
C8280 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 3.55e-19
C8281 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 9.94e-21
C8282 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 6.56e-21
C8283 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 5.84e-21
C8284 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# -8.41e-19
C8285 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 1.86e-21
C8286 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 7.69e-20
C8287 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 1.98e-19
C8288 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/Q_N 1.98e-19
C8289 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# V_LOW -0.00196f
C8290 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_1672_329# 1.07e-21
C8291 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0161f
C8292 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# -1.89e-19
C8293 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 2.84e-32
C8294 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# -2.37e-19
C8295 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_16_2/Y 2.81e-21
C8296 sky130_fd_sc_hd__inv_1_107/Y sky130_fd_sc_hd__inv_1_108/Y 1.93e-19
C8297 RISING_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00445f
C8298 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_1_20/Y 1.61e-19
C8299 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# V_LOW 0.0204f
C8300 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# CLOCK_GEN.SR_Op.Q 4.24e-21
C8301 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__inv_1_13/Y -7.92e-20
C8302 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_46/HI 0.00545f
C8303 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# sky130_fd_sc_hd__conb_1_36/HI 1.49e-19
C8304 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__inv_1_8/Y 0.00648f
C8305 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# V_LOW 0.0101f
C8306 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# V_GND -0.022f
C8307 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 0.00402f
C8308 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 1.19e-19
C8309 sky130_fd_sc_hd__inv_1_112/Y sky130_fd_sc_hd__inv_1_58/Y 1.17e-19
C8310 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 3.01e-21
C8311 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 0.00464f
C8312 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__conb_1_34/HI 0.0024f
C8313 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.29e-19
C8314 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__inv_1_53/Y 8.77e-20
C8315 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# V_GND 1.9e-19
C8316 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__conb_1_41/HI -3.05e-20
C8317 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__inv_1_90/Y 1.82e-19
C8318 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_2/A 0.0377f
C8319 sky130_fd_sc_hd__conb_1_44/LO V_LOW 0.00437f
C8320 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 2.05e-21
C8321 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 2.44e-20
C8322 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 6.3e-19
C8323 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/Q_N -9.56e-20
C8324 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__conb_1_40/LO 4.61e-20
C8325 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0401f
C8326 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_94/Y 0.0053f
C8327 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00678f
C8328 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# V_GND 0.00199f
C8329 sky130_fd_sc_hd__dfbbn_1_6/a_891_329# sky130_fd_sc_hd__inv_1_15/Y 1.23e-19
C8330 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__conb_1_5/LO 8.84e-20
C8331 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__conb_1_2/LO 3.77e-20
C8332 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 7.91e-19
C8333 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0.00204f
C8334 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 0.00204f
C8335 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__conb_1_18/LO 0.00106f
C8336 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# V_GND 0.00332f
C8337 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_0/HI 0.00804f
C8338 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# sky130_fd_sc_hd__inv_1_15/Y 5.43e-20
C8339 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.163f
C8340 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 8.58e-19
C8341 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 0.0682f
C8342 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_16/Y 0.0653f
C8343 sky130_fd_sc_hd__inv_1_11/Y V_LOW 0.0162f
C8344 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/Q_N -2.17e-19
C8345 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__inv_1_103/Y 4.15e-22
C8346 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# V_GND 0.00232f
C8347 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__inv_1_108/Y 6.44e-19
C8348 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0199f
C8349 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.00129f
C8350 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_16/Y 7.88e-21
C8351 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# V_LOW 3.29e-20
C8352 sky130_fd_sc_hd__inv_1_78/A sky130_fd_sc_hd__inv_1_86/Y 4.74e-20
C8353 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_68/A 2.11e-19
C8354 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 9.56e-22
C8355 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.29e-20
C8356 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# -0.242f
C8357 sky130_fd_sc_hd__inv_1_17/Y V_GND 0.155f
C8358 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.54e-20
C8359 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 1.86e-20
C8360 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 3.11e-19
C8361 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 2.73e-21
C8362 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 1.2e-20
C8363 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 8.63e-20
C8364 sky130_fd_sc_hd__dfbbn_1_32/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00307f
C8365 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_35/HI 0.00307f
C8366 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 3.72e-20
C8367 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 2.23e-20
C8368 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 0.00466f
C8369 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00715f
C8370 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 7.39e-19
C8371 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 2.11e-20
C8372 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# -0.00141f
C8373 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00339f
C8374 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 6.68e-20
C8375 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.11e-19
C8376 FALLING_COUNTER.COUNT_SUB_DFF7.Q V_LOW 1.28f
C8377 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 5.74e-20
C8378 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# sky130_fd_sc_hd__inv_16_1/Y 7.55e-20
C8379 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0124f
C8380 sky130_fd_sc_hd__conb_1_22/HI V_LOW 0.198f
C8381 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__inv_1_23/Y 2.55e-21
C8382 sky130_fd_sc_hd__conb_1_40/HI V_GND 0.105f
C8383 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0306f
C8384 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# V_GND 3.44e-19
C8385 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__conb_1_51/HI 1.56e-20
C8386 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 9.72e-20
C8387 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 3.35e-20
C8388 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 1.92e-20
C8389 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 6.33e-20
C8390 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0.00122f
C8391 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.44e-20
C8392 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# 2.74e-21
C8393 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 7.16e-19
C8394 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# 1.81e-19
C8395 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__conb_1_33/LO 2.6e-19
C8396 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.0173f
C8397 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_36/LO 0.0535f
C8398 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF17.Q 0.219f
C8399 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 0.00157f
C8400 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0355f
C8401 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0282f
C8402 sky130_fd_sc_hd__conb_1_19/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00323f
C8403 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 8.52e-21
C8404 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.38e-19
C8405 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 4.07e-21
C8406 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 6.79e-21
C8407 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.41e-19
C8408 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 3.18e-20
C8409 sky130_fd_sc_hd__dfbbn_1_27/Q_N RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0301f
C8410 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__conb_1_46/HI 0.00107f
C8411 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__inv_1_80/A 1.32e-19
C8412 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__conb_1_2/HI 0.00214f
C8413 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# V_LOW 0.0142f
C8414 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0297f
C8415 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# -1.66e-19
C8416 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__inv_1_103/Y 2.65e-21
C8417 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# sky130_fd_sc_hd__inv_1_20/Y 1.85e-19
C8418 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 3.07e-19
C8419 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_47/LO 0.0101f
C8420 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_35/LO 2.07e-19
C8421 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# sky130_fd_sc_hd__inv_1_13/Y 4.49e-21
C8422 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_47/HI 0.00114f
C8423 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_15/Y 5.74e-19
C8424 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# V_LOW 1.79e-20
C8425 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 3.69e-20
C8426 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# V_GND 3.02e-19
C8427 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.27e-20
C8428 transmission_gate_0/GN V_HIGH 0.224f
C8429 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# 3.27e-19
C8430 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00389f
C8431 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_85/A 8.98e-21
C8432 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 1.62e-20
C8433 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 9.45e-22
C8434 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 0.00118f
C8435 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 2.81e-20
C8436 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# 7.6e-19
C8437 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 0.00136f
C8438 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 0.00339f
C8439 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.0062f
C8440 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_26/LO 8.84e-20
C8441 sky130_fd_sc_hd__nand2_8_2/a_27_47# V_LOW -0.0089f
C8442 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# V_LOW 0.0131f
C8443 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.24e-21
C8444 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 5.02e-19
C8445 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 2.62e-21
C8446 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 4.01e-19
C8447 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00102f
C8448 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__inv_1_17/Y 1.82e-20
C8449 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# sky130_fd_sc_hd__inv_16_1/Y 3.79e-19
C8450 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# V_GND -6.56e-19
C8451 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00414f
C8452 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# -0.00441f
C8453 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.00724f
C8454 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.16e-20
C8455 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_101/Y 0.182f
C8456 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 4e-19
C8457 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# 4e-19
C8458 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# 5.51e-19
C8459 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# V_GND 3.2e-19
C8460 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00222f
C8461 sky130_fd_sc_hd__inv_2_0/Y V_GND 1.36f
C8462 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 1.81e-19
C8463 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 0.00207f
C8464 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 0.00443f
C8465 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 1.81e-19
C8466 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 0.00443f
C8467 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__conb_1_9/LO 0.00126f
C8468 sky130_fd_sc_hd__dfbbn_1_13/Q_N V_GND -0.00522f
C8469 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__inv_1_108/Y 4.54e-19
C8470 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# V_GND -0.00104f
C8471 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__conb_1_22/HI 0.00104f
C8472 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# V_GND 0.00643f
C8473 sky130_fd_sc_hd__inv_1_93/Y sky130_fd_sc_hd__inv_1_95/Y 5.55e-20
C8474 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 4.06e-21
C8475 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# sky130_fd_sc_hd__inv_1_47/Y 0.0112f
C8476 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# 9.85e-19
C8477 sky130_fd_sc_hd__inv_1_85/A V_GND 0.0866f
C8478 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# V_GND 0.00763f
C8479 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 4.55e-20
C8480 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__conb_1_45/HI 3.05e-21
C8481 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# sky130_fd_sc_hd__inv_16_1/Y 1.43e-20
C8482 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 4.07e-20
C8483 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 3.42e-20
C8484 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.34e-19
C8485 sky130_fd_sc_hd__conb_1_26/LO sky130_fd_sc_hd__inv_16_0/Y 0.00193f
C8486 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00142f
C8487 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__conb_1_0/HI 0.00326f
C8488 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# V_GND 0.00823f
C8489 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00214f
C8490 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_473_413# 4.05e-21
C8491 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00286f
C8492 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__dfbbn_1_5/a_581_47# 9.07e-21
C8493 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0353f
C8494 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__conb_1_51/HI 5.33e-21
C8495 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 3.87e-19
C8496 sky130_fd_sc_hd__inv_1_65/Y sky130_fd_sc_hd__inv_16_2/Y 1.76e-19
C8497 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.06e-20
C8498 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.249f
C8499 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 1.68e-19
C8500 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF9.Q 5.46e-20
C8501 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.00411f
C8502 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_23/Y 5.25e-21
C8503 sky130_fd_sc_hd__conb_1_50/HI V_LOW 0.193f
C8504 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.00571f
C8505 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 9.99e-20
C8506 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.86e-21
C8507 sky130_fd_sc_hd__fill_4_74/VPB V_GND 0.42f
C8508 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.613f
C8509 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__conb_1_33/HI 1.22e-20
C8510 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# sky130_fd_sc_hd__conb_1_2/HI 5.39e-19
C8511 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# -2.53e-20
C8512 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 1.61e-19
C8513 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_61/Y 9.32e-20
C8514 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__inv_1_20/Y 0.00648f
C8515 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_70/Y 0.214f
C8516 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__inv_1_15/Y 6.31e-21
C8517 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# V_GND 3.83e-19
C8518 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.336f
C8519 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.09e-20
C8520 sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 2.77e-20
C8521 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00141f
C8522 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 4.75e-21
C8523 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 1.43e-21
C8524 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# 5.21e-19
C8525 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.69e-20
C8526 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__conb_1_45/HI 2.13e-19
C8527 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.27e-21
C8528 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0661f
C8529 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# V_LOW 2.26e-20
C8530 sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__inv_1_70/A 9.07e-20
C8531 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# V_LOW -0.00389f
C8532 sky130_fd_sc_hd__inv_1_70/Y V_GND 0.081f
C8533 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.33e-19
C8534 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_17/Y 0.0236f
C8535 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_75/A 2.84e-20
C8536 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 2.63e-19
C8537 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 6.62e-21
C8538 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.45e-20
C8539 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# V_LOW 1.38e-19
C8540 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 7.69e-21
C8541 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# -3.03e-19
C8542 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# -0.00199f
C8543 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__inv_1_100/Y 0.00544f
C8544 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00312f
C8545 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__conb_1_0/HI 2.67e-20
C8546 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 0.003f
C8547 sky130_fd_sc_hd__dfbbn_1_45/a_891_329# V_LOW -0.00121f
C8548 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 5.01e-19
C8549 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__conb_1_22/LO 0.0179f
C8550 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_86/Y 0.0209f
C8551 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 6.04e-19
C8552 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.01e-20
C8553 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# -1.44e-20
C8554 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# 0.00215f
C8555 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.17e-19
C8556 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 0.549f
C8557 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__inv_16_2/Y 4.36e-20
C8558 sky130_fd_sc_hd__conb_1_11/HI sky130_fd_sc_hd__conb_1_12/HI 0.00118f
C8559 sky130_fd_sc_hd__dfbbn_1_18/a_891_329# V_LOW 2.26e-20
C8560 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__inv_1_119/Y 5.25e-19
C8561 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__inv_1_76/A 0.00639f
C8562 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# V_GND 5.73e-19
C8563 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# V_GND -0.00447f
C8564 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# V_LOW 0.00727f
C8565 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__conb_1_28/LO 1.35e-20
C8566 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_891_329# -2.2e-20
C8567 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# -3.48e-20
C8568 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# 0.00614f
C8569 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# V_GND 0.0066f
C8570 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_18/HI 0.0204f
C8571 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# V_GND 7.66e-19
C8572 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 6.8e-21
C8573 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_97/Y 0.0951f
C8574 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# V_GND 0.00172f
C8575 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -7.6e-19
C8576 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# -2.14e-19
C8577 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# V_LOW 0.0103f
C8578 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0.00111f
C8579 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00206f
C8580 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00144f
C8581 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# -5.54e-21
C8582 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# -9.62e-19
C8583 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -7.6e-19
C8584 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_381_47# 0.0187f
C8585 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# V_GND -0.00447f
C8586 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 4.28e-19
C8587 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_9/Y 1.67e-20
C8588 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__inv_1_59/Y 0.00417f
C8589 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# V_GND 4.02e-19
C8590 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0356f
C8591 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.00181f
C8592 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__conb_1_42/HI 1.1e-20
C8593 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# Reset 2.81e-19
C8594 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 8.85e-20
C8595 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 7.15e-19
C8596 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.134f
C8597 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_21/a_193_47# 8.09e-19
C8598 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 0.00787f
C8599 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__conb_1_24/HI 6.8e-19
C8600 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# V_LOW 2.26e-20
C8601 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# V_GND 0.00333f
C8602 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 0.00168f
C8603 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# -0.00122f
C8604 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# -0.00901f
C8605 sky130_fd_sc_hd__conb_1_17/LO FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0189f
C8606 sky130_fd_sc_hd__dfbbn_1_4/Q_N FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0273f
C8607 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.00326f
C8608 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.11e-19
C8609 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__dfbbn_1_39/Q_N 4.31e-20
C8610 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_1_108/Y 4.77e-20
C8611 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0121f
C8612 sky130_fd_sc_hd__dfbbn_1_29/a_1363_47# sky130_fd_sc_hd__conb_1_33/HI 1.35e-19
C8613 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.343f
C8614 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.75e-20
C8615 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# -1.44e-20
C8616 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__nand3_1_1/Y 0.0136f
C8617 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.44e-19
C8618 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -6.23e-21
C8619 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_381_47# -4.37e-20
C8620 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_42/a_941_21# -9.88e-20
C8621 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 4.43e-21
C8622 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 1.31e-19
C8623 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0011f
C8624 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_75/A 0.00308f
C8625 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__inv_1_62/Y 0.0159f
C8626 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1112_329# -0.00336f
C8627 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_381_47# -3.79e-20
C8628 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__inv_1_60/Y 0.00139f
C8629 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# V_GND 0.00171f
C8630 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__inv_1_11/Y 0.00943f
C8631 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__inv_16_0/Y 2.55e-19
C8632 FULL_COUNTER.COUNT_SUB_DFF4.Q V_LOW 1.1f
C8633 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/Q_N 7.36e-19
C8634 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 8.81e-20
C8635 sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# sky130_fd_sc_hd__inv_1_17/Y 5.83e-19
C8636 sky130_fd_sc_hd__nand2_8_5/a_27_47# V_LOW -0.00778f
C8637 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0199f
C8638 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_13/HI 0.0684f
C8639 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# V_LOW 0.0216f
C8640 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0435f
C8641 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.17e-19
C8642 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# V_LOW -0.00389f
C8643 FULL_COUNTER.COUNT_SUB_DFF7.Q V_LOW 1.23f
C8644 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 7.27e-20
C8645 sky130_fd_sc_hd__dfbbn_1_51/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.38e-19
C8646 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0015f
C8647 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 0.00123f
C8648 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# 0.00123f
C8649 sky130_fd_sc_hd__conb_1_25/LO RISING_COUNTER.COUNT_SUB_DFF4.Q 1.59e-19
C8650 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__conb_1_25/HI 0.0031f
C8651 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0174f
C8652 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# sky130_fd_sc_hd__inv_1_17/Y 7.97e-21
C8653 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.34e-19
C8654 FALLING_COUNTER.COUNT_SUB_DFF15.Q V_GND 1.66f
C8655 sky130_fd_sc_hd__inv_1_31/Y V_SENSE 0.0472f
C8656 sky130_fd_sc_hd__dfbbn_1_35/a_891_329# sky130_fd_sc_hd__inv_1_105/Y 6.1e-21
C8657 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.4e-20
C8658 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 1.42e-32
C8659 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# -0.00142f
C8660 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.89e-20
C8661 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# V_GND -0.00156f
C8662 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 0.00326f
C8663 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__conb_1_17/HI 4.43e-21
C8664 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_1_11/Y 8.88e-20
C8665 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF1.Q 9.35e-20
C8666 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.0439f
C8667 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# V_LOW 0.0691f
C8668 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# -6.43e-20
C8669 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# -3.06e-20
C8670 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00185f
C8671 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# -9.32e-20
C8672 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_891_329# 5.6e-21
C8673 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# V_GND 6.85e-19
C8674 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0443f
C8675 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 1.1e-19
C8676 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0.00502f
C8677 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0885f
C8678 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF15.Q 5.06e-20
C8679 sky130_fd_sc_hd__dfbbn_1_2/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.22e-19
C8680 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# -9.32e-20
C8681 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_941_21# -5.6e-19
C8682 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_473_413# -0.0103f
C8683 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.325f
C8684 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 4.03e-21
C8685 sky130_fd_sc_hd__conb_1_5/HI V_GND 0.133f
C8686 sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0266f
C8687 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0403f
C8688 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 0.0022f
C8689 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 4.55e-22
C8690 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# Reset 4.57e-19
C8691 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 3.07e-19
C8692 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.64e-19
C8693 sky130_fd_sc_hd__dfbbn_1_4/Q_N FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00418f
C8694 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.035f
C8695 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 9.16e-20
C8696 sky130_fd_sc_hd__inv_1_43/A V_LOW 0.342f
C8697 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0.00141f
C8698 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_21/a_193_47# 0.0104f
C8699 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# V_GND 0.00944f
C8700 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00287f
C8701 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# -3.79e-20
C8702 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# -0.00336f
C8703 sky130_fd_sc_hd__dfbbn_1_0/Q_N sky130_fd_sc_hd__inv_1_18/Y 2.73e-20
C8704 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# 2.49e-19
C8705 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# V_GND 0.00202f
C8706 RISING_COUNTER.COUNT_SUB_DFF2.Q V_GND 1.04f
C8707 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__conb_1_20/HI 0.00685f
C8708 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 3.29e-19
C8709 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0264f
C8710 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 1.77e-20
C8711 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.46e-20
C8712 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# -2.37e-19
C8713 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# -5.77e-20
C8714 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 2.84e-32
C8715 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_891_329# 8.64e-19
C8716 Reset FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.48e-21
C8717 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_60/Y 0.0875f
C8718 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_93/A 0.0019f
C8719 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__conb_1_30/HI 8.28e-19
C8720 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 0.00572f
C8721 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_59/Y 0.00165f
C8722 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__conb_1_4/LO 0.0144f
C8723 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 7.06e-19
C8724 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_557_413# -3.67e-20
C8725 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# -5.33e-20
C8726 sky130_fd_sc_hd__inv_1_78/A V_GND 0.153f
C8727 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0.00693f
C8728 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 2.28e-19
C8729 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# -4.66e-20
C8730 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# -3.79e-20
C8731 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0212f
C8732 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.11e-20
C8733 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_473_413# 0.00101f
C8734 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_381_47# -3.79e-20
C8735 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# -0.00336f
C8736 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00489f
C8737 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# V_LOW -1.01e-19
C8738 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.0023f
C8739 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 3.99e-19
C8740 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/Q_N -9.56e-20
C8741 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.042f
C8742 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 4.3e-20
C8743 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 3.31e-21
C8744 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__inv_1_4/Y 0.0484f
C8745 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 5.18e-21
C8746 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 4.81e-21
C8747 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 2.34e-21
C8748 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 7.84e-22
C8749 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__nand2_1_3/Y 9.37e-20
C8750 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 3.69e-20
C8751 sky130_fd_sc_hd__dfbbn_1_43/a_557_413# sky130_fd_sc_hd__inv_1_90/Y 8.17e-19
C8752 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00118f
C8753 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.46e-19
C8754 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__inv_1_9/Y 1.57e-20
C8755 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# V_GND 0.00501f
C8756 sky130_fd_sc_hd__dfbbn_1_44/Q_N V_LOW 2.15e-19
C8757 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 8.92e-19
C8758 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# V_GND 6.75e-19
C8759 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 3.89e-20
C8760 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.085f
C8761 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# sky130_fd_sc_hd__inv_16_2/Y 8.95e-19
C8762 sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# V_LOW 2.94e-20
C8763 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 5.99e-21
C8764 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__conb_1_41/HI 0.00104f
C8765 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 0.0335f
C8766 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/Q_N -4.24e-20
C8767 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.045f
C8768 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_106/Y 6.57e-20
C8769 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0.11f
C8770 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q -1.71e-20
C8771 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0.00145f
C8772 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.53e-19
C8773 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0537f
C8774 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 3.95e-20
C8775 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 1.8e-20
C8776 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/Q_N -4.33e-20
C8777 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.0417f
C8778 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# -6.8e-19
C8779 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 4.97e-19
C8780 sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0285f
C8781 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.6e-20
C8782 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_99/Y 0.15f
C8783 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.54e-20
C8784 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# sky130_fd_sc_hd__inv_1_19/Y 4.04e-19
C8785 sky130_fd_sc_hd__dfbbn_1_10/Q_N FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0242f
C8786 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_92/Y 0.00143f
C8787 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0198f
C8788 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 3.48e-21
C8789 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# V_GND 7.41e-19
C8790 FULL_COUNTER.COUNT_SUB_DFF14.Q V_GND 4.75f
C8791 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__conb_1_30/LO 2.82e-21
C8792 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__conb_1_28/HI 1.73e-19
C8793 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# sky130_fd_sc_hd__conb_1_20/HI 0.00115f
C8794 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00239f
C8795 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.00359f
C8796 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_42/HI 0.00226f
C8797 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 2.06e-20
C8798 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 1.09e-20
C8799 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 2.56e-20
C8800 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.92e-20
C8801 sky130_fd_sc_hd__nand3_1_2/a_109_47# sky130_fd_sc_hd__nand3_1_2/B 4.9e-19
C8802 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_101/Y 0.00745f
C8803 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# -1.66e-19
C8804 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 4.71e-20
C8805 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_557_413# 1.44e-19
C8806 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# 1.17e-19
C8807 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 4.61e-20
C8808 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 6.03e-20
C8809 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 6.53e-20
C8810 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# -1.63e-19
C8811 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__conb_1_8/HI 0.00315f
C8812 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 7.41e-21
C8813 sky130_fd_sc_hd__conb_1_18/LO FULL_COUNTER.COUNT_SUB_DFF8.Q 0.03f
C8814 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 9.19e-22
C8815 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0066f
C8816 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.85e-19
C8817 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 1.39e-20
C8818 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_76/A 0.0866f
C8819 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 7.61e-20
C8820 sky130_fd_sc_hd__dfbbn_1_39/a_891_329# V_LOW -0.00121f
C8821 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_83/Y 0.0329f
C8822 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__inv_1_53/Y 0.00333f
C8823 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.17e-20
C8824 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_12/Y 4.06e-21
C8825 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_11/HI 5.4e-19
C8826 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.029f
C8827 sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 9.39e-19
C8828 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# sky130_fd_sc_hd__conb_1_6/HI 0.00386f
C8829 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__conb_1_8/HI 3.29e-19
C8830 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00296f
C8831 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 1.02e-20
C8832 sky130_fd_sc_hd__inv_16_0/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 2.13e-20
C8833 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# 4.02e-19
C8834 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.2e-19
C8835 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# CLOCK_GEN.SR_Op.Q 4.87e-21
C8836 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.05e-19
C8837 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# V_LOW -0.104f
C8838 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# CLOCK_GEN.SR_Op.Q 0.166f
C8839 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_1_21/Y 1.62e-19
C8840 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 3.56e-19
C8841 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_12/HI 0.00158f
C8842 sky130_fd_sc_hd__dfbbn_1_31/Q_N FALLING_COUNTER.COUNT_SUB_DFF4.Q 8.34e-21
C8843 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.00532f
C8844 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00169f
C8845 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# V_GND 0.00171f
C8846 sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__conb_1_35/HI 0.0248f
C8847 sky130_fd_sc_hd__dfbbn_1_27/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 3.2e-21
C8848 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.18e-19
C8849 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.35e-19
C8850 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00213f
C8851 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__conb_1_31/HI 5.38e-19
C8852 RISING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_30/HI 7.37e-20
C8853 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 3.52e-19
C8854 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 1.73e-19
C8855 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 0.0357f
C8856 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 9.04e-21
C8857 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.45e-19
C8858 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# sky130_fd_sc_hd__inv_1_106/Y 8.96e-21
C8859 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 9.98e-20
C8860 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0907f
C8861 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 0.0389f
C8862 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 5.02e-20
C8863 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0.00133f
C8864 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_17/HI 2.12e-20
C8865 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.32e-19
C8866 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_18/Y 0.16f
C8867 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0369f
C8868 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1_22/LO 1.55e-20
C8869 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00379f
C8870 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# V_GND 0.00409f
C8871 Reset sky130_fd_sc_hd__inv_1_97/A 0.00318f
C8872 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.584f
C8873 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_1_112/Y 6.01e-21
C8874 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_75/A 6.27e-19
C8875 FULL_COUNTER.COUNT_SUB_DFF19.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0894f
C8876 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0353f
C8877 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__inv_1_102/Y 1.54e-19
C8878 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 0.00621f
C8879 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__conb_1_27/HI 1.37e-19
C8880 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_94/A 0.0895f
C8881 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00351f
C8882 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 0.0314f
C8883 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__conb_1_28/HI 2.03e-20
C8884 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0.00187f
C8885 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__conb_1_51/LO 0.00277f
C8886 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 9.04e-19
C8887 sky130_fd_sc_hd__inv_1_95/Y V_GND 0.0323f
C8888 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__inv_1_23/Y 0.236f
C8889 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 1.23e-19
C8890 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 9.28e-19
C8891 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# -1.61e-20
C8892 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_473_413# -3.86e-20
C8893 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 6.47e-19
C8894 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.072f
C8895 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__inv_1_98/Y 0.04f
C8896 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_16_0/Y 0.0188f
C8897 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_80/A 5.89e-20
C8898 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_16_1/Y 3.06e-19
C8899 RISING_COUNTER.COUNT_SUB_DFF3.Q V_LOW 3.52f
C8900 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0152f
C8901 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.82e-19
C8902 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 8.14e-20
C8903 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 1.52e-19
C8904 sky130_fd_sc_hd__inv_1_3/A V_GND 1.52f
C8905 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# 1.23e-19
C8906 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00243f
C8907 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.49e-21
C8908 sky130_fd_sc_hd__conb_1_44/LO FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.51e-20
C8909 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 0.0189f
C8910 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 5.06e-20
C8911 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__nand3_1_2/B 5.14e-19
C8912 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0123f
C8913 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__conb_1_30/HI 0.00123f
C8914 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF7.Q 0.592f
C8915 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# -3.72e-19
C8916 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# -5.77e-20
C8917 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# V_LOW -2.68e-19
C8918 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# CLOCK_GEN.SR_Op.Q 0.00228f
C8919 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.43e-21
C8920 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.43e-20
C8921 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 4.31e-19
C8922 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 2.11e-19
C8923 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__dfbbn_1_46/Q_N 3.82e-20
C8924 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 8.76e-22
C8925 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 0.0213f
C8926 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__inv_1_100/Y 0.0588f
C8927 sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__inv_1_9/Y 7.52e-22
C8928 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__inv_16_2/Y 4.18e-19
C8929 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_22/HI 2.37e-20
C8930 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.199f
C8931 sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# sky130_fd_sc_hd__inv_1_54/Y 3.75e-21
C8932 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.77e-20
C8933 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__conb_1_39/HI 1.01e-19
C8934 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 3.45e-20
C8935 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__conb_1_39/LO 0.00126f
C8936 sky130_fd_sc_hd__fill_4_58/VPB V_LOW 0.797f
C8937 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.28e-20
C8938 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# V_LOW 0.00427f
C8939 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__nand2_8_9/Y 4.6e-20
C8940 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00495f
C8941 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__conb_1_26/HI 1.11e-20
C8942 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 6.22e-19
C8943 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# V_LOW 0.0299f
C8944 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_102/Y 1.81e-20
C8945 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_473_413# -0.012f
C8946 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -0.00932f
C8947 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.58e-19
C8948 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# V_GND 2.83e-19
C8949 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.6e-19
C8950 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00289f
C8951 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0553f
C8952 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 0.00543f
C8953 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 4.21e-20
C8954 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__conb_1_28/HI 0.00126f
C8955 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 6.77e-20
C8956 sky130_fd_sc_hd__inv_1_4/Y V_LOW 0.332f
C8957 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 0.624f
C8958 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_57/Y 0.0275f
C8959 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# V_LOW 0.014f
C8960 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# 2.09e-19
C8961 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# V_GND 0.0022f
C8962 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.0201f
C8963 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# V_GND 0.00866f
C8964 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.44e-20
C8965 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# V_LOW 0.00905f
C8966 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0015f
C8967 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 1.71e-19
C8968 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0313f
C8969 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_95/A 1.16e-20
C8970 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# V_LOW 0.00694f
C8971 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# V_GND 0.00995f
C8972 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.14e-21
C8973 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# sky130_fd_sc_hd__conb_1_21/HI 3.23e-20
C8974 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 5.39e-19
C8975 RISING_COUNTER.COUNT_SUB_DFF13.Q V_LOW 1.08f
C8976 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_40/HI 0.0378f
C8977 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 9.29e-21
C8978 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 8.39e-20
C8979 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 1.56e-19
C8980 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# -3.79e-20
C8981 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# -0.00336f
C8982 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 2.84e-32
C8983 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI 5.85e-21
C8984 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# -2.57e-20
C8985 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__inv_1_6/Y 0.0107f
C8986 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 2.77e-20
C8987 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__inv_1_107/Y 5.67e-21
C8988 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00153f
C8989 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 4.14e-19
C8990 sky130_fd_sc_hd__dfbbn_1_33/a_581_47# sky130_fd_sc_hd__inv_1_98/Y 3.73e-19
C8991 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# V_GND 3.41e-19
C8992 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_70/A 0.00164f
C8993 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__inv_1_56/Y 0.0105f
C8994 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.31e-19
C8995 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# V_GND 0.00187f
C8996 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# V_LOW 0.038f
C8997 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0297f
C8998 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.67e-21
C8999 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# V_GND 0.00562f
C9000 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 9.53e-19
C9001 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# V_LOW 0.0048f
C9002 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 2.09e-20
C9003 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00102f
C9004 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 6.23e-22
C9005 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 9.54e-21
C9006 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# 0.00519f
C9007 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__conb_1_28/HI -1.31e-19
C9008 sky130_fd_sc_hd__conb_1_26/LO V_GND -0.00478f
C9009 FULL_COUNTER.COUNT_SUB_DFF1.Q V_GND 5.39f
C9010 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# -2.53e-20
C9011 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# -9.25e-19
C9012 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# -0.0103f
C9013 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__conb_1_26/HI 6.33e-19
C9014 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__inv_1_94/A 5.56e-19
C9015 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__conb_1_16/HI 8.48e-19
C9016 sky130_fd_sc_hd__inv_1_91/A V_LOW 0.146f
C9017 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 8.64e-20
C9018 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# sky130_fd_sc_hd__conb_1_30/HI -0.00125f
C9019 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 2.58e-20
C9020 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# -1.66e-19
C9021 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 5.14e-19
C9022 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -1.61e-19
C9023 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# -0.00834f
C9024 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_2/A 0.0223f
C9025 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/Y 0.33f
C9026 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# V_LOW 0.00299f
C9027 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_891_329# 0.00207f
C9028 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# V_GND -0.00397f
C9029 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 5.22e-19
C9030 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 2.62e-19
C9031 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# sky130_fd_sc_hd__conb_1_22/HI 4.94e-19
C9032 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# V_GND -0.00406f
C9033 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# -0.00813f
C9034 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# sky130_fd_sc_hd__conb_1_39/HI 2.71e-21
C9035 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__conb_1_38/HI 0.0116f
C9036 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.18e-20
C9037 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 3.61e-19
C9038 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 2.81e-19
C9039 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# V_LOW 1.74e-19
C9040 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.97e-19
C9041 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# V_LOW 2.26e-20
C9042 FALLING_COUNTER.COUNT_SUB_DFF14.Q V_GND 1.1f
C9043 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# V_LOW -6.55e-19
C9044 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# sky130_fd_sc_hd__inv_1_102/Y 5.14e-21
C9045 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 8.11e-21
C9046 FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_16_2/Y 0.124f
C9047 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1340_413# -2.57e-20
C9048 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_43/Y 2.06e-20
C9049 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.54e-19
C9050 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# V_GND -0.00806f
C9051 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.99e-19
C9052 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_88/Y 8.36e-20
C9053 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.12e-20
C9054 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0238f
C9055 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_39/HI -0.00236f
C9056 sky130_fd_sc_hd__dfbbn_1_50/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00383f
C9057 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 1.86e-21
C9058 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# CLOCK_GEN.SR_Op.Q 5.27e-19
C9059 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# 6.21e-20
C9060 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.68e-20
C9061 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 9.12e-21
C9062 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_97/A 2.61e-19
C9063 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_76/A 0.183f
C9064 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_1_18/Y 0.0144f
C9065 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 0.00152f
C9066 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_381_47# -2.53e-20
C9067 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_18/HI 4.17e-19
C9068 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# V_LOW 5.86e-19
C9069 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 0.0354f
C9070 sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# V_GND 1.59e-19
C9071 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00155f
C9072 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# V_GND 0.00179f
C9073 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# -0.00922f
C9074 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.11e-19
C9075 sky130_fd_sc_hd__dfbbn_1_0/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.06e-19
C9076 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__conb_1_35/HI 0.0137f
C9077 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# V_GND 6.86e-19
C9078 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__conb_1_24/LO 7.69e-20
C9079 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_54/Y 2.3e-20
C9080 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 2.73e-19
C9081 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 6.69e-20
C9082 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 2.07e-19
C9083 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 8.24e-19
C9084 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 8.33e-21
C9085 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__conb_1_0/HI 1.69e-20
C9086 sky130_fd_sc_hd__dfbbn_1_51/a_1340_413# sky130_fd_sc_hd__conb_1_40/HI 4.53e-19
C9087 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 8.14e-20
C9088 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.2e-21
C9089 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.021f
C9090 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00703f
C9091 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 2.11e-22
C9092 sky130_fd_sc_hd__conb_1_40/HI sky130_fd_sc_hd__inv_1_100/Y 2.68e-20
C9093 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__conb_1_44/HI 2.19e-20
C9094 FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_1/Y 0.193f
C9095 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00936f
C9096 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.89e-21
C9097 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__inv_1_4/Y 2.97e-19
C9098 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# V_GND 0.00147f
C9099 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# V_LOW 2.94e-20
C9100 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# sky130_fd_sc_hd__conb_1_38/HI 0.00134f
C9101 sky130_fd_sc_hd__conb_1_2/LO V_LOW 0.0874f
C9102 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# V_GND 0.00339f
C9103 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# V_LOW -6.55e-19
C9104 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 1.17e-19
C9105 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# 3.09e-19
C9106 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 0.00183f
C9107 sky130_fd_sc_hd__inv_16_1/Y V_LOW 5.64f
C9108 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 5.18e-19
C9109 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# sky130_fd_sc_hd__conb_1_28/HI 4.32e-20
C9110 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.11e-21
C9111 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0642f
C9112 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# -1.44e-20
C9113 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# -6.8e-19
C9114 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_9/LO 0.0478f
C9115 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.07e-20
C9116 sky130_fd_sc_hd__inv_1_72/A V_GND 0.158f
C9117 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# sky130_fd_sc_hd__conb_1_16/HI 4.33e-19
C9118 sky130_fd_sc_hd__inv_1_14/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 9.18e-20
C9119 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI 1.65e-19
C9120 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__conb_1_26/HI 6.89e-20
C9121 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# -0.00798f
C9122 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__conb_1_17/HI 0.0429f
C9123 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# -2.57e-20
C9124 sky130_fd_sc_hd__conb_1_29/LO V_LOW 0.0599f
C9125 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 9.36e-19
C9126 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_41/LO 0.00582f
C9127 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.5e-21
C9128 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# V_GND -0.00151f
C9129 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__inv_16_1/Y 1.38e-19
C9130 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.95e-19
C9131 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# V_GND -0.00157f
C9132 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# -1.44e-20
C9133 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_50/Y 0.111f
C9134 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# V_LOW -0.0167f
C9135 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_193_47# -1.71e-20
C9136 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# V_LOW 0.013f
C9137 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_31/HI 0.0384f
C9138 sky130_fd_sc_hd__conb_1_47/LO sky130_fd_sc_hd__inv_16_1/Y 2.34e-19
C9139 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__conb_1_17/HI 1.72e-20
C9140 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# -0.00144f
C9141 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# 0.00364f
C9142 sky130_fd_sc_hd__dfbbn_1_30/a_891_329# sky130_fd_sc_hd__conb_1_40/HI 9.76e-19
C9143 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 5.29e-21
C9144 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 0.0877f
C9145 sky130_fd_sc_hd__conb_1_19/HI V_LOW 0.166f
C9146 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# V_GND -0.0112f
C9147 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0303f
C9148 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0944f
C9149 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__conb_1_16/HI 0.00159f
C9150 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 5.22e-20
C9151 sky130_fd_sc_hd__conb_1_28/LO V_GND 0.00288f
C9152 sky130_fd_sc_hd__conb_1_4/HI V_GND 0.0456f
C9153 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 1.83e-20
C9154 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/Q_N 4.97e-19
C9155 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 9.8e-19
C9156 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 5.82e-20
C9157 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__inv_1_18/Y 6.87e-19
C9158 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.41e-21
C9159 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.19e-19
C9160 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# 0.00104f
C9161 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# -1.44e-20
C9162 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__inv_1_76/A 0.0117f
C9163 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.46e-19
C9164 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# V_GND 0.00575f
C9165 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# V_GND -0.00159f
C9166 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_16/HI 4.21e-21
C9167 sky130_fd_sc_hd__conb_1_39/LO V_GND 0.0033f
C9168 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_581_47# -2.6e-20
C9169 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# V_LOW 0.0134f
C9170 sky130_fd_sc_hd__dfbbn_1_22/a_891_329# sky130_fd_sc_hd__conb_1_32/HI 0.00119f
C9171 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.7e-19
C9172 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__conb_1_35/HI 0.00144f
C9173 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_36/HI 0.0976f
C9174 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_112/Y 0.0305f
C9175 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.324f
C9176 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# -3.79e-20
C9177 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1112_329# -0.00336f
C9178 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 2.44e-21
C9179 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 7.65e-21
C9180 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00112f
C9181 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 2.8e-20
C9182 sky130_fd_sc_hd__inv_1_83/Y V_LOW 0.528f
C9183 sky130_fd_sc_hd__nand2_8_6/a_27_47# Reset 0.00451f
C9184 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_107/Y 0.16f
C9185 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__inv_1_5/Y 1.67e-19
C9186 sky130_fd_sc_hd__dfbbn_1_11/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.9e-19
C9187 sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0235f
C9188 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 9.87e-21
C9189 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_1_58/Y 1.31e-20
C9190 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -5.77e-20
C9191 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# -2.37e-19
C9192 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 2.84e-32
C9193 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_112/Y 0.422f
C9194 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_65/Y 7.44e-19
C9195 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand2_8_9/Y 0.456f
C9196 sky130_fd_sc_hd__dfbbn_1_38/Q_N V_GND 0.00263f
C9197 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# V_GND -0.00934f
C9198 sky130_fd_sc_hd__dfbbn_1_50/Q_N V_GND 0.00182f
C9199 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# 0.00807f
C9200 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_2/Y 0.19f
C9201 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__inv_1_9/Y 5e-19
C9202 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__inv_16_0/Y 0.0364f
C9203 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.41e-19
C9204 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 5.55e-21
C9205 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0144f
C9206 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 5.67e-20
C9207 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 0.0192f
C9208 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_99/Y 0.00427f
C9209 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# sky130_fd_sc_hd__inv_1_63/Y 2.2e-19
C9210 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_193_47# -0.17f
C9211 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__conb_1_34/LO 9.15e-20
C9212 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__conb_1_44/HI 8.83e-20
C9213 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.13e-19
C9214 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# CLOCK_GEN.SR_Op.Q 2.68e-19
C9215 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_581_47# -7.91e-19
C9216 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 2.01e-19
C9217 sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# sky130_fd_sc_hd__conb_1_17/HI 4.8e-19
C9218 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_26/HI 0.0853f
C9219 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.02e-19
C9220 sky130_fd_sc_hd__conb_1_34/HI V_LOW 0.188f
C9221 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_67/Y 8.92e-20
C9222 sky130_fd_sc_hd__inv_1_40/A sky130_fd_sc_hd__inv_1_45/A 0.00134f
C9223 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 7.65e-20
C9224 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 3.75e-19
C9225 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__conb_1_48/HI 0.0128f
C9226 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# sky130_fd_sc_hd__inv_1_55/Y 7.1e-19
C9227 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# V_LOW -0.00522f
C9228 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# -3.72e-21
C9229 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# -0.0103f
C9230 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__conb_1_46/LO 9.17e-19
C9231 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.85e-21
C9232 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 7.89e-20
C9233 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# V_LOW -1.01e-19
C9234 sky130_fd_sc_hd__inv_1_108/Y V_GND 0.235f
C9235 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# -0.00107f
C9236 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__inv_1_57/Y 3.86e-19
C9237 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.85e-19
C9238 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_26/LO 3.72e-20
C9239 sky130_fd_sc_hd__conb_1_31/LO V_LOW 0.0485f
C9240 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 9.78e-20
C9241 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__conb_1_16/HI 2.03e-19
C9242 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_76/A 1.32f
C9243 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0302f
C9244 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__conb_1_28/HI 0.00222f
C9245 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 9.12e-19
C9246 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00124f
C9247 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 2.04e-19
C9248 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 6.62e-21
C9249 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__conb_1_26/HI 2.46e-20
C9250 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_1_102/Y 1.74e-19
C9251 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_74/Y 7.67e-20
C9252 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 0.00436f
C9253 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# V_LOW 0.0153f
C9254 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.61e-20
C9255 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_72/Y 0.157f
C9256 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# sky130_fd_sc_hd__inv_1_100/Y 5.99e-21
C9257 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0151f
C9258 sky130_fd_sc_hd__conb_1_4/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 5.02e-21
C9259 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/Q_N 8.52e-20
C9260 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# V_GND 0.00944f
C9261 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# 0.00619f
C9262 sky130_fd_sc_hd__conb_1_42/LO V_LOW 0.0953f
C9263 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 2.46e-19
C9264 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_20/LO 0.0367f
C9265 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 3.67e-19
C9266 sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# V_GND 6.32e-19
C9267 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# V_GND -0.0135f
C9268 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0611f
C9269 CLOCK_GEN.SR_Op.Q Reset 0.709f
C9270 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__nor2_1_0/Y 1.8e-20
C9271 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.46e-20
C9272 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# 0.0366f
C9273 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 3.6e-20
C9274 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 3.63e-20
C9275 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# sky130_fd_sc_hd__inv_1_112/Y 0.00222f
C9276 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__inv_1_107/Y 0.0368f
C9277 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__conb_1_32/LO 1.28e-19
C9278 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# sky130_fd_sc_hd__nand3_1_2/Y 8.26e-19
C9279 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00145f
C9280 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_40/HI 0.0259f
C9281 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_93/A 0.104f
C9282 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_19/HI 8.06e-21
C9283 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 1.79e-21
C9284 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__conb_1_0/HI 0.0323f
C9285 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# V_GND -0.0473f
C9286 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_36/HI 0.00674f
C9287 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__inv_1_103/Y 0.00568f
C9288 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# -1.66e-19
C9289 sky130_fd_sc_hd__nand2_8_8/a_27_47# Reset 0.242f
C9290 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.419f
C9291 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# Reset 1.5e-19
C9292 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_1_100/Y 1.66e-20
C9293 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__inv_1_61/Y 0.00318f
C9294 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# CLOCK_GEN.SR_Op.Q 4.06e-21
C9295 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# V_GND -0.0135f
C9296 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__conb_1_34/HI 0.00633f
C9297 sky130_fd_sc_hd__conb_1_11/LO sky130_fd_sc_hd__conb_1_11/HI 0.00486f
C9298 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 6.05e-20
C9299 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_42/HI 0.0192f
C9300 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0111f
C9301 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 6.79e-21
C9302 sky130_fd_sc_hd__conb_1_37/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 8.16e-19
C9303 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# -0.00385f
C9304 sky130_fd_sc_hd__conb_1_1/LO V_GND -0.00353f
C9305 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__inv_1_59/Y 5.86e-19
C9306 sky130_fd_sc_hd__dfbbn_1_20/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0207f
C9307 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__conb_1_9/LO 7.33e-21
C9308 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# 6.66e-20
C9309 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__conb_1_24/HI -6.47e-19
C9310 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 2.58e-20
C9311 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00628f
C9312 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00109f
C9313 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.0214f
C9314 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__conb_1_37/HI 2.46e-19
C9315 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_2/HI 0.00649f
C9316 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# -0.0242f
C9317 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 1.15e-19
C9318 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 0.00193f
C9319 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__conb_1_48/HI 0.0238f
C9320 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__inv_1_4/Y 0.0049f
C9321 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_22/Y 2.47e-21
C9322 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0226f
C9323 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__conb_1_41/HI 8.56e-22
C9324 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 4.85e-21
C9325 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 8.86e-22
C9326 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# V_LOW -6.55e-19
C9327 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0579f
C9328 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_51/A 7.11e-20
C9329 sky130_fd_sc_hd__inv_1_3/Y V_GND 0.02f
C9330 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# sky130_fd_sc_hd__conb_1_5/HI 0.00144f
C9331 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 2.02e-20
C9332 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_791_47# 3.23e-20
C9333 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# V_LOW -0.0013f
C9334 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# 2.05e-19
C9335 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__inv_1_98/Y 1.66e-19
C9336 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_96/A 0.0181f
C9337 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 1.31e-22
C9338 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_57/Y 0.0253f
C9339 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 5.96e-19
C9340 sky130_fd_sc_hd__dfbbn_1_16/a_1112_329# sky130_fd_sc_hd__conb_1_4/HI 0.00306f
C9341 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.12f
C9342 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 1.45e-22
C9343 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.0059f
C9344 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 1.32e-19
C9345 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 6.03e-19
C9346 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 1.78e-19
C9347 sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# V_GND 0.00126f
C9348 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 3.02e-20
C9349 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00549f
C9350 FULL_COUNTER.COUNT_SUB_DFF2.Q V_GND 6.98f
C9351 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# 0.00399f
C9352 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 1.19e-20
C9353 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 7.39e-21
C9354 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 0.00658f
C9355 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.0305f
C9356 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.0194f
C9357 FALLING_COUNTER.COUNT_SUB_DFF0.Q V_LOW 1.23f
C9358 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_10/HI -0.00233f
C9359 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00303f
C9360 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# 2.97e-19
C9361 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# V_GND 3.01e-19
C9362 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# -0.0323f
C9363 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_10/HI 0.00405f
C9364 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 9.06e-19
C9365 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# V_GND 2.81e-19
C9366 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 9.54e-20
C9367 sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# sky130_fd_sc_hd__conb_1_36/HI 5.75e-19
C9368 sky130_fd_sc_hd__dfbbn_1_37/a_581_47# sky130_fd_sc_hd__inv_1_103/Y 0.00108f
C9369 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_24/LO 0.00869f
C9370 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# Reset 3.37e-19
C9371 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 2.29e-22
C9372 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.562f
C9373 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# sky130_fd_sc_hd__inv_1_61/Y 1.07e-21
C9374 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__conb_1_34/LO 4.5e-21
C9375 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__conb_1_11/HI 5.28e-20
C9376 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__inv_1_100/Y 3.97e-20
C9377 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_59/Y 0.0101f
C9378 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# sky130_fd_sc_hd__conb_1_34/HI 8.88e-20
C9379 sky130_fd_sc_hd__conb_1_13/HI V_LOW 0.0265f
C9380 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00195f
C9381 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# sky130_fd_sc_hd__conb_1_42/HI 9.74e-19
C9382 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# V_GND -0.176f
C9383 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_23/LO 0.00131f
C9384 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_17/HI 0.00424f
C9385 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__conb_1_24/HI 0.00264f
C9386 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 0.0357f
C9387 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.52e-21
C9388 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 8.27e-21
C9389 sky130_fd_sc_hd__conb_1_36/LO V_LOW 0.0761f
C9390 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 0.0012f
C9391 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 1.67e-21
C9392 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__inv_1_56/Y 0.0124f
C9393 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_1_11/Y 0.0131f
C9394 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.61e-19
C9395 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# V_GND 0.0449f
C9396 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.45e-21
C9397 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# sky130_fd_sc_hd__inv_1_108/Y 1.64e-19
C9398 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00262f
C9399 sky130_fd_sc_hd__conb_1_47/LO V_LOW 0.0951f
C9400 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_45/Q_N 0.0242f
C9401 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__inv_1_21/Y 0.041f
C9402 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 1.26e-20
C9403 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 2.65e-20
C9404 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_1_105/Y 4.24e-20
C9405 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0463f
C9406 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.00617f
C9407 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 8.05e-20
C9408 sky130_fd_sc_hd__conb_1_29/HI V_GND 0.107f
C9409 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.84e-19
C9410 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# -0.0182f
C9411 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.63e-20
C9412 sky130_fd_sc_hd__conb_1_51/HI sky130_fd_sc_hd__conb_1_38/HI 2.07e-20
C9413 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_891_329# 7.75e-19
C9414 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.77e-21
C9415 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# sky130_fd_sc_hd__conb_1_5/HI 3.52e-19
C9416 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.81e-19
C9417 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_22/HI 1.47e-19
C9418 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00584f
C9419 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 2.24e-20
C9420 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__conb_1_42/HI 8.45e-19
C9421 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__conb_1_30/HI 1.66e-20
C9422 Reset sky130_fd_sc_hd__inv_1_97/Y 0.00132f
C9423 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0313f
C9424 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 3.32e-20
C9425 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_68/A 1.2e-19
C9426 sky130_fd_sc_hd__inv_1_119/Y sky130_fd_sc_hd__inv_2_0/Y 2.07f
C9427 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0.0106f
C9428 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0145f
C9429 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# V_GND -0.154f
C9430 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_94/A 1.44e-19
C9431 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_941_21# -0.0014f
C9432 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# -2.37e-19
C9433 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__inv_1_22/Y 0.00337f
C9434 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00188f
C9435 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# V_LOW 0.00647f
C9436 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# V_LOW 0.0223f
C9437 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_1/LO 0.00223f
C9438 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/Q_N 0.0249f
C9439 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__conb_1_27/HI 0.00116f
C9440 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_9/Y 0.245f
C9441 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__inv_1_105/Y 9.07e-19
C9442 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00107f
C9443 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# 1.45e-19
C9444 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 0.00212f
C9445 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 3.89e-19
C9446 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.4e-21
C9447 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_60/Y 0.0669f
C9448 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# V_LOW -8.74e-19
C9449 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__nand2_8_9/Y 1.99e-19
C9450 sky130_fd_sc_hd__dfbbn_1_3/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.52e-19
C9451 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# V_LOW -9.15e-19
C9452 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# sky130_fd_sc_hd__conb_1_9/HI -0.00741f
C9453 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__conb_1_10/HI 1.51e-19
C9454 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_68/A 1.56e-19
C9455 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_19/LO 8.59e-21
C9456 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_20/Y 1.2e-19
C9457 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_70/A 0.0123f
C9458 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__conb_1_47/HI 0.0161f
C9459 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_24/LO 0.00169f
C9460 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# 0.0104f
C9461 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_891_329# 3.56e-21
C9462 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.46e-19
C9463 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__conb_1_14/LO 1.31e-20
C9464 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_48/LO 7.32e-19
C9465 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# sky130_fd_sc_hd__conb_1_11/HI -6.57e-19
C9466 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# V_LOW 3.56e-20
C9467 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# V_GND 9.32e-19
C9468 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# -2.32e-19
C9469 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# -2.66e-19
C9470 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# V_LOW -0.0185f
C9471 sky130_fd_sc_hd__dfbbn_1_48/Q_N sky130_fd_sc_hd__conb_1_34/HI 1.17e-19
C9472 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# V_GND 0.00471f
C9473 sky130_fd_sc_hd__inv_1_21/Y V_GND 0.0805f
C9474 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# V_LOW 1.38e-19
C9475 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 0.0222f
C9476 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 0.00286f
C9477 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__inv_1_58/Y 3.69e-19
C9478 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.00507f
C9479 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# V_GND 0.00435f
C9480 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# V_GND 1.92e-19
C9481 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__conb_1_13/HI 6.22e-19
C9482 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# sky130_fd_sc_hd__inv_1_10/Y 9.58e-19
C9483 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.85e-19
C9484 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_647_21# -6.43e-20
C9485 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_473_413# -0.00985f
C9486 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# V_LOW 0.0106f
C9487 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_41/HI 4.22e-19
C9488 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__inv_1_47/Y 7.11e-20
C9489 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_37/HI 0.00306f
C9490 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_8_2/A 7.14e-19
C9491 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 3.46e-21
C9492 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.02e-21
C9493 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF6.Q 2.33e-19
C9494 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# V_GND 0.0102f
C9495 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.01e-19
C9496 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 7.56e-19
C9497 sky130_fd_sc_hd__conb_1_18/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0137f
C9498 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 2.69e-19
C9499 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0.00813f
C9500 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 4.17e-19
C9501 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 2.9e-20
C9502 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 0.001f
C9503 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 0.0174f
C9504 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00644f
C9505 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# V_GND 2.05e-19
C9506 FULL_COUNTER.COUNT_SUB_DFF16.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00163f
C9507 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_16_2/Y 2.32e-19
C9508 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__inv_1_22/Y 0.0933f
C9509 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# V_LOW 0.0134f
C9510 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# V_GND 1.86e-19
C9511 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 9.81e-21
C9512 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# V_LOW 0.0236f
C9513 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# V_GND 0.00114f
C9514 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# sky130_fd_sc_hd__inv_1_21/Y 1.86e-19
C9515 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# V_LOW 1.02e-19
C9516 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0163f
C9517 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00256f
C9518 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_91/Y 0.413f
C9519 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 7.36e-19
C9520 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# V_LOW -9.15e-19
C9521 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.62e-20
C9522 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# V_GND -0.0115f
C9523 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_27/HI 0.249f
C9524 FULL_COUNTER.COUNT_SUB_DFF18.Q V_GND 0.971f
C9525 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.15e-19
C9526 FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_41/HI 6.7e-20
C9527 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__conb_1_35/LO 1.29e-19
C9528 sky130_fd_sc_hd__inv_1_56/Y CLOCK_GEN.SR_Op.Q 3.46e-21
C9529 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 4.56e-20
C9530 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.25e-20
C9531 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 0.0298f
C9532 sky130_fd_sc_hd__inv_1_69/Y Reset 0.00292f
C9533 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# Reset 0.016f
C9534 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_1_62/Y 6.39e-21
C9535 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__inv_1_18/Y 0.0139f
C9536 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0.00108f
C9537 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 9.54e-19
C9538 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 4.99e-19
C9539 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 8.58e-21
C9540 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 1.43e-21
C9541 sky130_fd_sc_hd__dfbbn_1_10/Q_N V_LOW -0.0104f
C9542 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# V_GND -0.0474f
C9543 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 0.0306f
C9544 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__inv_1_76/A 9.17e-20
C9545 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# V_GND 0.00575f
C9546 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 0.00339f
C9547 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 3.59e-21
C9548 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# -5.72e-19
C9549 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# -0.0103f
C9550 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# V_GND -0.0038f
C9551 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 2.66e-19
C9552 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# V_LOW -0.322f
C9553 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# V_GND 1.15e-19
C9554 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# -1.66e-19
C9555 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# -5.16e-20
C9556 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__inv_1_58/Y 0.00716f
C9557 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0309f
C9558 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# V_LOW -1.39e-35
C9559 sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# V_LOW 2.94e-20
C9560 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_12/HI 0.0106f
C9561 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 1.91e-21
C9562 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0547f
C9563 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# sky130_fd_sc_hd__conb_1_27/HI 0.00196f
C9564 sky130_fd_sc_hd__dfbbn_1_34/Q_N sky130_fd_sc_hd__inv_1_105/Y 0.0104f
C9565 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 7.03e-19
C9566 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 2.84e-32
C9567 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# -2.52e-19
C9568 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -0.00164f
C9569 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__inv_1_75/A 4.85e-21
C9570 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_94/Y 1.55e-19
C9571 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/Q_N 5.15e-21
C9572 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 0.00163f
C9573 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 0.00949f
C9574 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.00949f
C9575 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 7.67e-19
C9576 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0.00163f
C9577 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 7.67e-19
C9578 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# sky130_fd_sc_hd__conb_1_9/HI -5.54e-19
C9579 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# V_LOW -9.15e-19
C9580 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 4.5e-19
C9581 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# V_LOW 0.00114f
C9582 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# sky130_fd_sc_hd__conb_1_47/HI 9.42e-19
C9583 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_647_21# -5.67e-19
C9584 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# V_GND -0.0141f
C9585 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# 0.04f
C9586 sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 8.3e-20
C9587 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__inv_1_12/Y 0.0025f
C9588 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__conb_1_13/HI 2.61e-19
C9589 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# -1.66e-19
C9590 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# -7.17e-20
C9591 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# V_LOW -0.0103f
C9592 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__inv_1_12/Y 0.0224f
C9593 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# V_GND 8.02e-19
C9594 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 0.0342f
C9595 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_891_329# -0.00159f
C9596 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# -0.00486f
C9597 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.13e-19
C9598 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_8/Y 4.06e-21
C9599 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 5.45e-21
C9600 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0179f
C9601 RISING_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00211f
C9602 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# 5.06e-19
C9603 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# V_GND 0.00578f
C9604 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0.358f
C9605 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_21/HI 8.85e-19
C9606 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_9/Y 0.00197f
C9607 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# sky130_fd_sc_hd__conb_1_13/HI -5.17e-19
C9608 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 6.48e-20
C9609 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# -0.00375f
C9610 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 3.03e-19
C9611 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/Q_N 1.59e-21
C9612 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_32/HI 0.0323f
C9613 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# V_GND 9.9e-20
C9614 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 7.94e-20
C9615 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# V_LOW -0.32f
C9616 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_21/HI 1.46e-19
C9617 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# V_GND -0.00273f
C9618 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.98e-20
C9619 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# sky130_fd_sc_hd__conb_1_34/HI 8.42e-19
C9620 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 2.53e-19
C9621 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 2.21e-21
C9622 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/Q_N 9.65e-21
C9623 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 2.6e-20
C9624 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_13/HI 8.96e-20
C9625 sky130_fd_sc_hd__dfbbn_1_48/a_581_47# Reset 3e-21
C9626 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_647_21# -1.27e-19
C9627 sky130_fd_sc_hd__nand2_1_0/a_113_47# Reset 5.15e-19
C9628 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_381_47# 2.11e-20
C9629 sky130_fd_sc_hd__conb_1_36/HI FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.117f
C9630 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__inv_1_103/Y 0.0437f
C9631 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00267f
C9632 sky130_fd_sc_hd__dfbbn_1_36/Q_N sky130_fd_sc_hd__inv_1_105/Y 0.00813f
C9633 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.2e-20
C9634 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_50/A 3.18e-19
C9635 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00282f
C9636 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 8.85e-20
C9637 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# V_GND -2.37e-19
C9638 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.0015f
C9639 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0.00158f
C9640 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.13e-19
C9641 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# V_GND 3.78e-19
C9642 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# Reset 0.0139f
C9643 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 4.97e-22
C9644 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.16e-22
C9645 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_16/HI 0.134f
C9646 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# V_GND -0.0458f
C9647 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__conb_1_41/HI 1.01e-19
C9648 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.0189f
C9649 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# -4.66e-20
C9650 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_381_47# -3.79e-20
C9651 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# Reset 1.91e-19
C9652 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 1.16e-19
C9653 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# V_GND 2.7e-19
C9654 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0917f
C9655 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00109f
C9656 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# V_GND 0.00564f
C9657 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.01f
C9658 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# -6.8e-19
C9659 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# -0.00119f
C9660 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# V_GND -0.00443f
C9661 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_22/HI 0.00218f
C9662 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# -1.03e-19
C9663 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_473_413# -3.86e-20
C9664 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 9.12e-19
C9665 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 2.04e-19
C9666 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 6.62e-21
C9667 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 0.00124f
C9668 V_GND V_SENSE 40.8f
C9669 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_97/Y 0.00727f
C9670 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_90/Y 1.01e-19
C9671 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_80/A 7.23e-20
C9672 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 0.00212f
C9673 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0.00212f
C9674 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# -0.0158f
C9675 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -6.4e-19
C9676 sky130_fd_sc_hd__dfbbn_1_48/Q_N V_LOW -0.00503f
C9677 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00357f
C9678 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 6.95e-20
C9679 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_23/LO 1.67e-19
C9680 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# -7.17e-20
C9681 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# -1.76e-19
C9682 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# -0.00151f
C9683 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# -2.32e-19
C9684 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 5.48e-21
C9685 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.76e-21
C9686 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# sky130_fd_sc_hd__inv_1_20/Y 3e-20
C9687 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.00501f
C9688 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 5.36e-19
C9689 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00501f
C9690 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 5.36e-19
C9691 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 1.72e-20
C9692 sky130_fd_sc_hd__dfbbn_1_18/Q_N sky130_fd_sc_hd__conb_1_9/HI -2.17e-19
C9693 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 7.4e-20
C9694 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__conb_1_44/HI 5.57e-19
C9695 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__conb_1_47/HI 3.29e-20
C9696 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 5.44e-21
C9697 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_86/Y 0.0262f
C9698 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# V_GND 2.14e-19
C9699 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__conb_1_2/HI 0.00372f
C9700 sky130_fd_sc_hd__dfbbn_1_12/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 3.77e-19
C9701 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__conb_1_22/HI 5.71e-21
C9702 sky130_fd_sc_hd__inv_1_16/Y V_LOW 0.0344f
C9703 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# sky130_fd_sc_hd__inv_1_12/Y 7.93e-19
C9704 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# 3.23e-21
C9705 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 6.31e-21
C9706 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 1.4e-21
C9707 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 8.95e-21
C9708 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__inv_1_12/Y 0.00109f
C9709 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.1e-20
C9710 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.61e-19
C9711 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# V_LOW -0.0863f
C9712 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# -3.46e-20
C9713 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 1.42e-32
C9714 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 5.74e-19
C9715 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__conb_1_39/HI 0.00115f
C9716 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_94/A 0.0139f
C9717 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0125f
C9718 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# V_LOW 4.8e-20
C9719 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# 3.13e-19
C9720 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.98e-20
C9721 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# sky130_fd_sc_hd__inv_1_9/Y 1.25e-19
C9722 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_41/HI 0.0584f
C9723 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_16_1/Y 0.399f
C9724 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# -0.00107f
C9725 sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# sky130_fd_sc_hd__conb_1_32/HI 1.57e-19
C9726 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0188f
C9727 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_68/A 0.00716f
C9728 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__nand2_8_9/Y 5.41e-19
C9729 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# V_GND -0.00357f
C9730 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 0.00368f
C9731 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 1.26e-21
C9732 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__conb_1_13/HI 5.5e-21
C9733 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 4.69e-20
C9734 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_15/Y 0.175f
C9735 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 9.61e-21
C9736 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 1.05e-19
C9737 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__conb_1_19/LO 0.0144f
C9738 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_581_47# -2.6e-20
C9739 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.1f
C9740 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# -2.65e-20
C9741 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 9.46e-22
C9742 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.55e-19
C9743 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# V_GND 0.00425f
C9744 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_97/A 0.0446f
C9745 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_12/LO 0.0164f
C9746 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# -0.00934f
C9747 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_0/A 0.613f
C9748 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# V_LOW 0.0232f
C9749 sky130_fd_sc_hd__dfbbn_1_1/Q_N FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00161f
C9750 sky130_fd_sc_hd__conb_1_39/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0333f
C9751 sky130_fd_sc_hd__dfbbn_1_46/a_581_47# V_GND -9.19e-19
C9752 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 6.48e-20
C9753 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 7.18e-20
C9754 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.45e-19
C9755 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 1.14e-21
C9756 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.15e-19
C9757 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.454f
C9758 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.72e-20
C9759 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# V_GND 3.34e-19
C9760 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__conb_1_41/HI 1.69e-19
C9761 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_68/A 0.00395f
C9762 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_581_47# 2.2e-19
C9763 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# -0.0189f
C9764 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_557_413# -0.0012f
C9765 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1_68/A 0.0451f
C9766 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 3.33e-19
C9767 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 2.93e-20
C9768 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 6.21e-20
C9769 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 7.69e-19
C9770 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 7.21e-19
C9771 sky130_fd_sc_hd__dfbbn_1_43/a_581_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.99e-19
C9772 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_8/Y 0.0291f
C9773 sky130_fd_sc_hd__conb_1_31/HI V_GND 0.551f
C9774 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_17/HI 1.12e-20
C9775 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_581_47# -2.6e-20
C9776 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# V_GND -0.0063f
C9777 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# sky130_fd_sc_hd__conb_1_51/HI 3.11e-19
C9778 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# -2.57e-20
C9779 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__inv_1_112/Y 0.109f
C9780 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_557_413# 1.93e-19
C9781 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__inv_1_76/A 1.47e-20
C9782 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_16/a_891_329# 1.72e-20
C9783 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 2.02e-20
C9784 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_791_47# 3.23e-20
C9785 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# V_LOW 0.0213f
C9786 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_891_329# 0.00292f
C9787 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__inv_1_12/Y 0.0061f
C9788 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 2.23e-19
C9789 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_1_53/Y 1.28e-20
C9790 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# -6.8e-19
C9791 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 3.49e-20
C9792 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 3.49e-20
C9793 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_105/Y 5.9e-19
C9794 sky130_fd_sc_hd__conb_1_32/HI sky130_fd_sc_hd__inv_16_1/Y 1.14e-20
C9795 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__nand3_1_2/B 0.182f
C9796 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 8.13e-20
C9797 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 0.00116f
C9798 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 3.43e-20
C9799 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 1.09e-20
C9800 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 4.45e-22
C9801 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# -7.17e-20
C9802 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# -1.64e-19
C9803 sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__inv_1_75/A 4.58e-21
C9804 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 8.26e-21
C9805 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# V_LOW -0.00294f
C9806 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 1.76e-19
C9807 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/Q_N 1.76e-19
C9808 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 7.65e-19
C9809 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 7.65e-19
C9810 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0023f
C9811 sky130_fd_sc_hd__inv_1_2/A V_SENSE 0.047f
C9812 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# -1.6e-19
C9813 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# -5.54e-21
C9814 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_1_20/Y 3.52e-19
C9815 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__conb_1_49/HI 0.0157f
C9816 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# V_LOW 9.32e-19
C9817 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# CLOCK_GEN.SR_Op.Q 1.57e-22
C9818 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__inv_1_8/Y 0.00373f
C9819 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__inv_1_13/Y 4.34e-20
C9820 sky130_fd_sc_hd__conb_1_44/LO FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0134f
C9821 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# sky130_fd_sc_hd__conb_1_22/HI 1.35e-21
C9822 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# V_GND 0.00812f
C9823 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# V_LOW 0.0205f
C9824 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 2.55e-19
C9825 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_50/Y 6.95e-20
C9826 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_71/A 6.62e-20
C9827 CLOCK_GEN.SR_Op.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 1e-19
C9828 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_557_413# 3.84e-19
C9829 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.45e-20
C9830 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# V_LOW -2.68e-19
C9831 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.8e-19
C9832 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__inv_1_53/Y 1.68e-19
C9833 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# V_GND 3.38e-19
C9834 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__inv_1_90/Y 7.72e-20
C9835 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 5.84e-19
C9836 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 0.00498f
C9837 sky130_fd_sc_hd__dfbbn_1_49/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00167f
C9838 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.00255f
C9839 sky130_fd_sc_hd__dfbbn_1_9/Q_N V_GND -0.00659f
C9840 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# V_GND 0.00393f
C9841 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__conb_1_5/LO 8.84e-20
C9842 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__conb_1_6/HI 2.54e-19
C9843 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 9.82e-20
C9844 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 5.61e-19
C9845 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# V_GND 4.16e-19
C9846 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0952f
C9847 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.00742f
C9848 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 0.00447f
C9849 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_16/Y 0.0263f
C9850 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# V_GND 8.91e-20
C9851 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__inv_1_108/Y 0.0107f
C9852 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__inv_1_16/Y 1.01e-19
C9853 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_581_47# -7.91e-19
C9854 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 1.05e-19
C9855 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 2.25e-19
C9856 sky130_fd_sc_hd__conb_1_50/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0103f
C9857 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_11/Y 3.37e-21
C9858 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# -0.0079f
C9859 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__conb_1_25/HI 9.82e-20
C9860 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0.00447f
C9861 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.69e-20
C9862 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 9.87e-19
C9863 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 0.00108f
C9864 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.00139f
C9865 sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 4.53e-19
C9866 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_35/HI 0.00113f
C9867 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0.00427f
C9868 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__conb_1_41/HI 9.45e-19
C9869 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 6.16e-19
C9870 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__conb_1_45/HI 7.15e-20
C9871 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 1.88e-19
C9872 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_1_20/Y 4.03e-19
C9873 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.0016f
C9874 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 1.92e-19
C9875 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.02e-21
C9876 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# sky130_fd_sc_hd__inv_16_1/Y 6.97e-19
C9877 sky130_fd_sc_hd__inv_1_62/Y RISING_COUNTER.COUNT_SUB_DFF9.Q 0.227f
C9878 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0431f
C9879 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__inv_1_23/Y 1.31e-20
C9880 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.76e-21
C9881 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 9.61e-20
C9882 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0143f
C9883 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# V_GND -0.0121f
C9884 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# sky130_fd_sc_hd__conb_1_34/HI 6.33e-20
C9885 sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# sky130_fd_sc_hd__conb_1_51/HI -2.65e-20
C9886 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 7.01e-21
C9887 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.47e-20
C9888 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 4.1e-20
C9889 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 1.09e-19
C9890 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0.0124f
C9891 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0.00799f
C9892 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 6.02e-19
C9893 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.204f
C9894 sky130_fd_sc_hd__dfbbn_1_13/a_1363_47# sky130_fd_sc_hd__inv_1_12/Y 4.63e-20
C9895 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.014f
C9896 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# 4.36e-21
C9897 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 3.32e-20
C9898 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 0.00628f
C9899 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 0.00766f
C9900 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0144f
C9901 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00694f
C9902 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_76/A 0.11f
C9903 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00184f
C9904 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 5.88e-20
C9905 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 3.17e-21
C9906 sky130_fd_sc_hd__conb_1_33/HI V_LOW 0.0304f
C9907 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.67e-19
C9908 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__conb_1_46/HI -0.00171f
C9909 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# V_LOW 5.39e-19
C9910 sky130_fd_sc_hd__inv_1_80/A V_LOW 0.45f
C9911 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__conb_1_2/HI 0.00525f
C9912 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.166f
C9913 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# -9.32e-20
C9914 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 1.49e-19
C9915 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# sky130_fd_sc_hd__conb_1_49/HI 0.00435f
C9916 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__conb_1_35/LO 9e-21
C9917 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__inv_1_103/Y 0.305f
C9918 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# sky130_fd_sc_hd__inv_1_8/Y 1.07e-21
C9919 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_47/HI 0.00577f
C9920 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__inv_1_15/Y 1.85e-21
C9921 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# V_GND 0.00562f
C9922 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# V_LOW 0.00145f
C9923 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__inv_1_100/Y 0.0132f
C9924 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.18e-20
C9925 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_1_57/Y 1.53e-20
C9926 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00402f
C9927 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00135f
C9928 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_381_47# 0.00455f
C9929 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 1.79e-19
C9930 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 1.97e-20
C9931 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 5.2e-20
C9932 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 1.29e-20
C9933 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 2.26e-20
C9934 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.79e-19
C9935 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__conb_1_39/HI 8.46e-20
C9936 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0362f
C9937 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__conb_1_45/HI 4.9e-19
C9938 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 7.65e-19
C9939 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 2.07e-19
C9940 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# V_LOW 0.00534f
C9941 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 4.1e-22
C9942 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__inv_1_53/Y 5.77e-19
C9943 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 7.11e-20
C9944 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 7.74e-19
C9945 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 1.73e-19
C9946 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.87e-19
C9947 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 0.00204f
C9948 sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__inv_16_0/Y 0.031f
C9949 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_2_0/Y 8.59e-19
C9950 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.231f
C9951 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# V_GND 0.00212f
C9952 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.00282f
C9953 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_891_329# -1.42e-19
C9954 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_557_413# -3.67e-20
C9955 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# -6.29e-19
C9956 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_1_54/Y 0.00218f
C9957 sky130_fd_sc_hd__conb_1_15/HI V_GND 0.0175f
C9958 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.048f
C9959 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 0.00162f
C9960 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 0.00102f
C9961 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 0.00521f
C9962 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 0.00521f
C9963 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 0.00102f
C9964 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 0.00162f
C9965 sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__nand2_1_0/Y 0.0595f
C9966 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# sky130_fd_sc_hd__inv_1_108/Y 8.91e-20
C9967 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# V_GND -0.00164f
C9968 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# V_GND -0.176f
C9969 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__conb_1_22/HI 0.00102f
C9970 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.0497f
C9971 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.158f
C9972 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_8/HI 0.00818f
C9973 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# V_GND 0.00367f
C9974 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# V_GND 0.0316f
C9975 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_581_47# -7.91e-19
C9976 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 3.12e-19
C9977 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 8.11e-21
C9978 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# 1.54e-19
C9979 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 2.02e-20
C9980 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.00188f
C9981 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# 8.11e-19
C9982 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# V_GND 0.00364f
C9983 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# sky130_fd_sc_hd__conb_1_35/HI 5.88e-20
C9984 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_97/A 0.00209f
C9985 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 1.81e-20
C9986 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 1.88e-19
C9987 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 8.11e-19
C9988 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 2.54e-20
C9989 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 4.5e-19
C9990 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 5.48e-19
C9991 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.82e-20
C9992 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__conb_1_0/HI 0.00108f
C9993 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# V_GND -3.91e-19
C9994 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 3.09e-19
C9995 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_941_21# 4.57e-20
C9996 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 1.94e-19
C9997 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0018f
C9998 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 6.27e-20
C9999 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand3_1_2/B 0.0145f
C10000 sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.21e-20
C10001 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00821f
C10002 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_99/Y 0.0861f
C10003 FALLING_COUNTER.COUNT_SUB_DFF5.Q V_GND 0.588f
C10004 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 3.47e-19
C10005 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 0.1f
C10006 sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.23e-20
C10007 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.347f
C10008 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__inv_16_2/Y 0.0468f
C10009 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_102/Y 0.00142f
C10010 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# 4.86e-21
C10011 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 3.13e-20
C10012 RISING_COUNTER.COUNT_SUB_DFF10.Q V_LOW 0.838f
C10013 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.00445f
C10014 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0258f
C10015 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00319f
C10016 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# sky130_fd_sc_hd__conb_1_46/HI 0.00142f
C10017 sky130_fd_sc_hd__dfbbn_1_5/Q_N V_LOW -0.00916f
C10018 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__conb_1_26/HI 8.84e-20
C10019 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# sky130_fd_sc_hd__conb_1_2/HI 1.1e-19
C10020 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00236f
C10021 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# -5.33e-20
C10022 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_557_413# -3.67e-20
C10023 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/Q_N -4.33e-20
C10024 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_21/Y 0.001f
C10025 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.561f
C10026 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__inv_1_20/Y 0.00373f
C10027 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 2.64e-21
C10028 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_104/Y 0.00218f
C10029 sky130_fd_sc_hd__inv_1_19/Y V_GND 0.048f
C10030 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# -0.0554f
C10031 sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0358f
C10032 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_95/A 0.00386f
C10033 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# V_GND 0.00339f
C10034 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__inv_1_11/Y 0.041f
C10035 FALLING_COUNTER.COUNT_SUB_DFF10.Q V_LOW 1.16f
C10036 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 5.29e-19
C10037 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00257f
C10038 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# 1.23e-19
C10039 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# 0.00104f
C10040 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# V_LOW 4.8e-20
C10041 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.97e-21
C10042 sky130_fd_sc_hd__dfbbn_1_26/a_557_413# V_LOW -9.15e-19
C10043 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.57e-19
C10044 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_891_329# 5.5e-20
C10045 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_17/Y 0.0244f
C10046 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 7.74e-21
C10047 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.13e-20
C10048 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# V_LOW 3.56e-20
C10049 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_381_47# -0.00375f
C10050 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_1_100/Y 3.36e-20
C10051 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00718f
C10052 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 0.00668f
C10053 sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# V_LOW -0.00266f
C10054 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_581_47# 5.35e-20
C10055 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 0.0014f
C10056 sky130_fd_sc_hd__dfbbn_1_43/Q_N V_GND -5.91e-19
C10057 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 4.01e-20
C10058 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# sky130_fd_sc_hd__inv_1_54/Y 1.15e-21
C10059 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00207f
C10060 FULL_COUNTER.COUNT_SUB_DFF16.Q V_LOW 1.4f
C10061 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 1.64e-19
C10062 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 9.29e-20
C10063 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_791_47# 2.17e-20
C10064 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 2.17e-20
C10065 sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# V_LOW 4.8e-20
C10066 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# V_GND -8.88e-19
C10067 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# V_GND 9.15e-20
C10068 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# V_LOW 1.38e-19
C10069 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_381_47# -3.79e-20
C10070 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# -4.66e-20
C10071 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# 0.00144f
C10072 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# V_GND 0.00179f
C10073 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_70/A 0.00406f
C10074 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# sky130_fd_sc_hd__conb_1_18/HI 1.69e-19
C10075 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_8/HI 1.44e-20
C10076 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# V_GND 1.68e-19
C10077 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__conb_1_28/HI 4.73e-22
C10078 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_50/Y 1.7e-20
C10079 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# V_GND 2.05e-19
C10080 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# V_LOW 0.00569f
C10081 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# V_GND 0.0182f
C10082 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# -6.22e-19
C10083 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# -6.23e-21
C10084 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# -0.00464f
C10085 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 4.82e-20
C10086 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.51e-19
C10087 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 2.02e-20
C10088 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 3.71e-20
C10089 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_381_47# -0.00464f
C10090 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# -1.67e-19
C10091 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__dfbbn_1_50/a_941_21# -6.22e-19
C10092 sky130_fd_sc_hd__inv_1_89/A V_GND 0.0139f
C10093 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_557_413# 4.94e-19
C10094 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# sky130_fd_sc_hd__conb_1_49/HI 1.71e-19
C10095 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 9.4e-21
C10096 sky130_fd_sc_hd__dfbbn_1_18/a_581_47# V_GND 2.65e-19
C10097 sky130_fd_sc_hd__conb_1_4/LO V_LOW 0.0943f
C10098 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1_46/HI 0.00443f
C10099 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0197f
C10100 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# V_GND 9.12e-19
C10101 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 1.32e-20
C10102 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# Reset 0.0112f
C10103 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.89e-19
C10104 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__inv_1_90/Y 6e-19
C10105 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.046f
C10106 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 7.34e-19
C10107 sky130_fd_sc_hd__conb_1_32/HI V_LOW 0.13f
C10108 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__conb_1_8/LO 0.00764f
C10109 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 0.00152f
C10110 sky130_fd_sc_hd__dfbbn_1_40/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 6.42e-19
C10111 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# -0.141f
C10112 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_16_1/Y 0.3f
C10113 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# V_LOW 4.8e-20
C10114 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# V_GND 0.00389f
C10115 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 1.04e-19
C10116 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_21/HI 1.33e-20
C10117 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_473_413# -0.00834f
C10118 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# -1.61e-19
C10119 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_45/A 0.0945f
C10120 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__inv_1_19/Y 6.39e-20
C10121 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.00116f
C10122 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00564f
C10123 sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00335f
C10124 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 6.59e-19
C10125 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.73e-19
C10126 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_76/A 8.67e-19
C10127 sky130_fd_sc_hd__conb_1_19/LO FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00577f
C10128 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 5.2e-19
C10129 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_10/Y 1.82e-19
C10130 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.34e-19
C10131 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.209f
C10132 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__inv_1_101/Y 0.00138f
C10133 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 8.84e-19
C10134 sky130_fd_sc_hd__dfbbn_1_1/Q_N sky130_fd_sc_hd__conb_1_2/HI 2.91e-19
C10135 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.39e-20
C10136 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 3.07e-21
C10137 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_381_47# -2.53e-20
C10138 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 8.86e-21
C10139 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__conb_1_40/HI 1.76e-19
C10140 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 9.64e-19
C10141 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# sky130_fd_sc_hd__inv_1_20/Y 1.07e-21
C10142 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_39/LO 2.03e-19
C10143 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 3.05e-21
C10144 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_16_1/Y 8.04e-20
C10145 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_54/Y 9.56e-20
C10146 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__inv_1_60/Y 2.33e-21
C10147 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# V_GND -9.15e-19
C10148 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# -0.134f
C10149 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_54/Y 3.48e-19
C10150 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.49e-19
C10151 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# sky130_fd_sc_hd__inv_1_17/Y 0.00255f
C10152 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0115f
C10153 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# V_LOW -0.312f
C10154 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# -0.179f
C10155 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.233f
C10156 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__conb_1_38/LO 1.53e-19
C10157 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_13/Y 2.21e-21
C10158 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# -0.00141f
C10159 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00365f
C10160 sky130_fd_sc_hd__dfbbn_1_19/a_557_413# V_LOW -9.15e-19
C10161 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# sky130_fd_sc_hd__inv_1_108/Y 1.4e-19
C10162 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_1_23/Y 0.4f
C10163 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_50/Q_N 4.01e-19
C10164 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.04e-20
C10165 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.51e-19
C10166 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 6.79e-20
C10167 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 1.16e-19
C10168 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.0136f
C10169 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# 5.33e-19
C10170 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 5.33e-19
C10171 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__conb_1_25/HI 4.62e-20
C10172 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00973f
C10173 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0311f
C10174 sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# sky130_fd_sc_hd__inv_1_105/Y 3.02e-21
C10175 sky130_fd_sc_hd__conb_1_40/LO FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0191f
C10176 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.16e-20
C10177 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.014f
C10178 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# V_GND -0.0405f
C10179 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_67/Y 3.79e-20
C10180 sky130_fd_sc_hd__dfbbn_1_15/Q_N V_GND 0.00208f
C10181 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__conb_1_18/HI 3e-19
C10182 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 9.25e-19
C10183 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_1_11/Y 0.00394f
C10184 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.0129f
C10185 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_25/HI 8.11e-21
C10186 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# V_LOW 0.0207f
C10187 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# -3.86e-20
C10188 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# -0.00341f
C10189 sky130_fd_sc_hd__conb_1_48/HI V_GND 0.451f
C10190 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.18e-19
C10191 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# 5.23e-21
C10192 sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# V_GND 1.13e-19
C10193 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0392f
C10194 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_74/Y 0.0257f
C10195 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__conb_1_49/HI 6.8e-19
C10196 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0179f
C10197 sky130_fd_sc_hd__conb_1_34/LO sky130_fd_sc_hd__conb_1_34/HI 0.0116f
C10198 sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__inv_1_119/Y 0.00546f
C10199 sky130_fd_sc_hd__dfbbn_1_2/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00121f
C10200 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_941_21# -0.00134f
C10201 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# -2.37e-19
C10202 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0392f
C10203 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_1_72/A 8.28e-20
C10204 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_1_106/Y 0.0182f
C10205 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00111f
C10206 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_19/Y 0.0974f
C10207 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 0.00256f
C10208 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# Reset 6.69e-19
C10209 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.46e-20
C10210 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 7.94e-20
C10211 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.1e-19
C10212 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 7.69e-20
C10213 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.71e-19
C10214 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0242f
C10215 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 1.16e-20
C10216 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# V_GND 0.0214f
C10217 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00626f
C10218 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# V_GND 0.0019f
C10219 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# -2.57e-20
C10220 sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__inv_1_1/Y 9.07e-20
C10221 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_3/Y 0.0229f
C10222 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 5.37e-22
C10223 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_23/LO 0.00154f
C10224 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_65/Y 1.31e-19
C10225 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_2_0/Y 8.28e-20
C10226 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.25e-19
C10227 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__conb_1_20/HI -0.054f
C10228 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0496f
C10229 sky130_fd_sc_hd__conb_1_51/HI FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.168f
C10230 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.55e-20
C10231 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0237f
C10232 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# -5.54e-21
C10233 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# 0.00389f
C10234 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# -1.44e-20
C10235 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_75/A 0.00247f
C10236 sky130_fd_sc_hd__conb_1_38/HI V_GND -0.179f
C10237 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_59/Y 3.31e-19
C10238 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# 0.00792f
C10239 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_891_329# -2.2e-20
C10240 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# -3.48e-20
C10241 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_17/LO 3.72e-20
C10242 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.69e-21
C10243 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 4.12e-19
C10244 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 4.78e-19
C10245 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_16_2/Y 0.109f
C10246 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_20/Y 0.0693f
C10247 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_18/Y 2.95e-19
C10248 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_75/Y 0.00966f
C10249 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 1.54e-19
C10250 sky130_fd_sc_hd__conb_1_42/LO sky130_fd_sc_hd__conb_1_45/LO 0.00297f
C10251 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.564f
C10252 sky130_fd_sc_hd__dfbbn_1_12/a_581_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.25e-19
C10253 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.132f
C10254 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 4.39e-19
C10255 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 1.29e-20
C10256 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__nand2_8_2/A 8.47e-21
C10257 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 2.24e-21
C10258 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 2.51e-19
C10259 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.63e-19
C10260 sky130_fd_sc_hd__conb_1_35/LO FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.83e-19
C10261 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.47e-22
C10262 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 2.22e-19
C10263 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 2.39e-21
C10264 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.97e-21
C10265 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# sky130_fd_sc_hd__inv_1_90/Y 7.05e-19
C10266 sky130_fd_sc_hd__dfbbn_1_21/a_1159_47# sky130_fd_sc_hd__conb_1_25/HI 0.00253f
C10267 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00367f
C10268 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__inv_1_9/Y 0.00419f
C10269 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00183f
C10270 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# V_GND 0.00462f
C10271 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_21/HI 4.56e-21
C10272 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00369f
C10273 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# V_GND 1.58e-19
C10274 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__inv_1_11/Y 0.0277f
C10275 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__conb_1_5/HI 8.83e-20
C10276 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 9.04e-19
C10277 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_50/Y 0.00692f
C10278 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_31/LO 0.0816f
C10279 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.57f
C10280 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# V_LOW 1.44e-19
C10281 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 6.52e-21
C10282 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# -2.57e-20
C10283 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__conb_1_37/HI 0.0115f
C10284 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/Q_N -9.56e-20
C10285 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.0417f
C10286 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q -3.39e-20
C10287 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__inv_1_106/Y 4.71e-20
C10288 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 0.0338f
C10289 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.49e-20
C10290 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00121f
C10291 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.00247f
C10292 sky130_fd_sc_hd__conb_1_12/HI V_GND -0.071f
C10293 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 3.29e-20
C10294 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 6e-19
C10295 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 4.54e-21
C10296 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.72e-19
C10297 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# -1.66e-19
C10298 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/Q_N -9.56e-20
C10299 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00112f
C10300 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_44/HI 0.0195f
C10301 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.00314f
C10302 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_42/Y 2.28e-19
C10303 RISING_COUNTER.COUNT_SUB_DFF11.Q CLOCK_GEN.SR_Op.Q 1.31e-20
C10304 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__nand3_1_0/Y 4.42e-20
C10305 sky130_fd_sc_hd__inv_1_99/Y V_LOW 0.247f
C10306 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.31e-20
C10307 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__conb_1_3/HI 4.6e-20
C10308 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 6.6e-19
C10309 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 4.67e-21
C10310 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.014f
C10311 sky130_fd_sc_hd__dfbbn_1_19/Q_N FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0255f
C10312 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_5/HI 1.65e-19
C10313 sky130_fd_sc_hd__inv_1_90/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0091f
C10314 RISING_COUNTER.COUNT_SUB_DFF5.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 8.17e-20
C10315 sky130_fd_sc_hd__inv_2_0/A V_GND 0.0813f
C10316 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 2.49e-19
C10317 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 1.09e-20
C10318 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 3.69e-19
C10319 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# V_GND 6.13e-19
C10320 sky130_fd_sc_hd__dfbbn_1_51/Q_N V_GND 0.00203f
C10321 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_95/A 2.8e-20
C10322 sky130_fd_sc_hd__nand2_1_5/Y V_GND 0.175f
C10323 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00398f
C10324 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__conb_1_28/HI 8.46e-21
C10325 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__inv_1_99/Y 0.00743f
C10326 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_1_60/Y 1.29e-19
C10327 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 8.42e-19
C10328 FULL_COUNTER.COUNT_SUB_DFF5.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 9.19e-20
C10329 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 3.49e-19
C10330 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_93/A 0.102f
C10331 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 2.54e-19
C10332 sky130_fd_sc_hd__dfbbn_1_24/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 7.64e-19
C10333 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF3.Q 6.05e-19
C10334 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.98e-20
C10335 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 1.02e-20
C10336 sky130_fd_sc_hd__nand3_1_2/a_193_47# sky130_fd_sc_hd__nand3_1_2/B 9.26e-19
C10337 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 8.51e-19
C10338 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 2.81f
C10339 sky130_fd_sc_hd__conb_1_18/HI V_GND 0.208f
C10340 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 4.57e-20
C10341 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 4.71e-19
C10342 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.37e-20
C10343 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.00109f
C10344 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 9.28e-19
C10345 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.00479f
C10346 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 1.42e-32
C10347 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# -3.46e-20
C10348 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.52e-20
C10349 sky130_fd_sc_hd__conb_1_49/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0314f
C10350 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.919f
C10351 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.56e-19
C10352 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_31/LO 3.11e-19
C10353 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 2.78e-19
C10354 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 1.34e-20
C10355 sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# V_LOW -0.00266f
C10356 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__inv_1_53/Y 1.81e-20
C10357 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0.00155f
C10358 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00249f
C10359 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 7.54e-19
C10360 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0512f
C10361 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.123f
C10362 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# sky130_fd_sc_hd__conb_1_6/HI 3.72e-19
C10363 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.44e-19
C10364 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_791_47# 3.78e-19
C10365 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0306f
C10366 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 2.37e-19
C10367 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 1.59e-20
C10368 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00114f
C10369 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand2_8_2/A 3.97e-19
C10370 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# CLOCK_GEN.SR_Op.Q 3.89e-20
C10371 sky130_fd_sc_hd__fill_4_63/VPB V_GND 0.437f
C10372 sky130_fd_sc_hd__conb_1_34/LO V_LOW 0.0915f
C10373 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF13.Q 3.82e-21
C10374 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.96e-19
C10375 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# V_LOW 0.00757f
C10376 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# CLOCK_GEN.SR_Op.Q 0.0735f
C10377 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_1_12/Y 0.117f
C10378 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 0.00174f
C10379 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__conb_1_12/HI 1.77e-19
C10380 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 4.35e-19
C10381 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00119f
C10382 sky130_fd_sc_hd__dfbbn_1_39/a_581_47# V_GND -9.04e-19
C10383 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_54/Y 0.0238f
C10384 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.83e-19
C10385 sky130_fd_sc_hd__conb_1_45/LO V_LOW 0.151f
C10386 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__conb_1_5/HI 3.64e-19
C10387 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 2.41e-19
C10388 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.00893f
C10389 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_97/Y 0.0484f
C10390 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_31/HI 1.03e-19
C10391 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__inv_1_11/Y 3.42e-19
C10392 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 4.1e-19
C10393 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__conb_1_26/HI 6.7e-19
C10394 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# sky130_fd_sc_hd__conb_1_37/HI 0.0174f
C10395 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 2.67e-20
C10396 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_63/Y 0.277f
C10397 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 6.23e-21
C10398 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.43e-20
C10399 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0266f
C10400 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_11/LO 3.64e-20
C10401 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 7.59e-20
C10402 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0355f
C10403 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 7.69e-20
C10404 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_18/Y 0.0926f
C10405 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 7.01e-21
C10406 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 1.48e-19
C10407 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# V_GND 1.92e-19
C10408 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 2.66e-19
C10409 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__conb_1_2/HI 1.36e-20
C10410 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0301f
C10411 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# sky130_fd_sc_hd__inv_1_108/Y 9.49e-20
C10412 sky130_fd_sc_hd__conb_1_43/HI V_LOW 0.209f
C10413 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__conb_1_42/HI 2.75e-19
C10414 sky130_fd_sc_hd__dfbbn_1_47/a_581_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00177f
C10415 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_63/Y 0.059f
C10416 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 0.0199f
C10417 FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_15/Y 0.046f
C10418 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.312f
C10419 sky130_fd_sc_hd__inv_1_94/Y V_LOW 0.484f
C10420 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.00164f
C10421 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_99/Y 8.05e-21
C10422 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 8.82e-20
C10423 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 0.0027f
C10424 sky130_fd_sc_hd__conb_1_9/HI V_GND -0.0816f
C10425 sky130_fd_sc_hd__dfbbn_1_15/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 1.12e-19
C10426 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 7.68e-20
C10427 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_46/LO 3.65e-20
C10428 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.00191f
C10429 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.00841f
C10430 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 3.86e-22
C10431 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_93/A 5.77e-20
C10432 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_75/A 0.0312f
C10433 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_16_1/Y 0.458f
C10434 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# -0.193f
C10435 RISING_COUNTER.COUNT_SUB_DFF8.Q V_LOW 3.3f
C10436 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# -2.37e-19
C10437 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_941_21# -3.01e-19
C10438 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 2.75e-21
C10439 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/Q_N -4.33e-20
C10440 sky130_fd_sc_hd__conb_1_0/HI V_LOW 0.161f
C10441 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0336f
C10442 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_51/A 8.34e-20
C10443 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/Q_N 0.00129f
C10444 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__inv_1_98/Y 0.0469f
C10445 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_42/HI 2.41e-21
C10446 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__inv_1_8/Y 4.88e-20
C10447 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 4.04e-19
C10448 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# sky130_fd_sc_hd__conb_1_34/LO 1.53e-19
C10449 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.99e-19
C10450 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__conb_1_28/LO 8.84e-20
C10451 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00445f
C10452 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 0.0373f
C10453 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_8_2/A 0.112f
C10454 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# 1.75e-19
C10455 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_2_0/Y 0.0421f
C10456 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_1/LO 8.84e-20
C10457 sky130_fd_sc_hd__conb_1_12/LO V_GND 6.51e-19
C10458 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00483f
C10459 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.25e-20
C10460 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0.162f
C10461 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__nand3_1_2/B 3.83e-19
C10462 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 2.17e-21
C10463 RISING_COUNTER.COUNT_SUB_DFF14.Q CLOCK_GEN.SR_Op.Q 4.33e-19
C10464 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__conb_1_30/HI -0.051f
C10465 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__inv_1_4/Y 3.93e-19
C10466 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# -2.01e-20
C10467 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# CLOCK_GEN.SR_Op.Q 8.69e-22
C10468 sky130_fd_sc_hd__inv_16_0/Y Reset 0.0724f
C10469 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# V_LOW -7.16e-19
C10470 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# CLOCK_GEN.SR_Op.Q 0.0184f
C10471 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.93e-20
C10472 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.85e-21
C10473 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 7.72e-22
C10474 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 1.88e-20
C10475 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 5.32e-19
C10476 sky130_fd_sc_hd__conb_1_8/LO FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00534f
C10477 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 3e-20
C10478 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_22/HI 0.387f
C10479 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 1.96e-19
C10480 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.63e-19
C10481 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_112/Y 5.65e-20
C10482 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0715f
C10483 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.04e-20
C10484 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.58e-20
C10485 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__conb_1_39/HI 1.48e-21
C10486 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__inv_1_9/Y 3.85e-19
C10487 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 8.12e-19
C10488 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 9.78e-19
C10489 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 7.19e-19
C10490 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__nand2_8_9/Y 1.4e-19
C10491 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# V_LOW 0.0204f
C10492 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__conb_1_31/HI 8.52e-21
C10493 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00795f
C10494 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__conb_1_26/HI 3.48e-20
C10495 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__conb_1_37/HI 0.0301f
C10496 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 2.77e-20
C10497 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__conb_1_6/HI 1.39e-20
C10498 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# V_LOW -0.312f
C10499 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0139f
C10500 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0321f
C10501 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/Q_N 0.0231f
C10502 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_102/Y 2.29e-19
C10503 sky130_fd_sc_hd__dfbbn_1_29/Q_N RISING_COUNTER.COUNT_SUB_DFF2.Q 6.99e-20
C10504 sky130_fd_sc_hd__dfbbn_1_40/Q_N FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0284f
C10505 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# -2.52e-19
C10506 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -0.0114f
C10507 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 2.49e-19
C10508 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# sky130_fd_sc_hd__inv_1_18/Y 7.59e-19
C10509 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 6.69e-19
C10510 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 4.47e-20
C10511 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0779f
C10512 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 5.48e-21
C10513 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__nand2_8_3/Y 0.0148f
C10514 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 4.68e-21
C10515 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 3.2e-19
C10516 sky130_fd_sc_hd__inv_1_91/Y Reset 0.582f
C10517 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF0.Q 0.473f
C10518 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# V_LOW 0.00315f
C10519 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_57/Y 0.0278f
C10520 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# 3.98e-19
C10521 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# V_GND 3.03e-19
C10522 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_51/Y 4.94e-19
C10523 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 0.014f
C10524 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF19.Q 2.55e-19
C10525 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00199f
C10526 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# V_GND 0.0106f
C10527 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# V_LOW 0.0119f
C10528 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.54e-19
C10529 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.37f
C10530 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0306f
C10531 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_23/Y 1.83e-20
C10532 sky130_fd_sc_hd__inv_1_62/Y V_GND 0.0143f
C10533 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_22/Y 0.00779f
C10534 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_16_2/Y 0.276f
C10535 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_14/LO 4.91e-19
C10536 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# V_LOW -0.0376f
C10537 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# V_GND 0.00422f
C10538 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00164f
C10539 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__conb_1_21/HI 3.66e-19
C10540 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_40/HI 0.0328f
C10541 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.00165f
C10542 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 9.97e-20
C10543 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 5.65e-19
C10544 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 9.96e-19
C10545 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_71/Y 1.69e-19
C10546 sky130_fd_sc_hd__conb_1_0/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0787f
C10547 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__conb_1_30/HI 0.00132f
C10548 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# -1.66e-19
C10549 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF19.Q 0.00148f
C10550 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.73e-21
C10551 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# sky130_fd_sc_hd__inv_1_6/Y 3.12e-19
C10552 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_1_107/Y 2.29e-21
C10553 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_43/A 2.78e-19
C10554 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_17/HI 3.53e-20
C10555 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00373f
C10556 sky130_fd_sc_hd__conb_1_29/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 4.79e-19
C10557 FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_16_2/Y 0.111f
C10558 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__inv_1_59/Y 3.01e-19
C10559 sky130_fd_sc_hd__conb_1_6/LO V_LOW 0.0924f
C10560 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# V_GND 4.61e-19
C10561 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_41/HI 0.0335f
C10562 sky130_fd_sc_hd__inv_1_54/Y V_LOW 0.202f
C10563 sky130_fd_sc_hd__inv_1_0/A V_SENSE 0.0667f
C10564 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# V_GND 0.00181f
C10565 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.49e-20
C10566 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# V_LOW 0.00875f
C10567 sky130_fd_sc_hd__dfbbn_1_14/Q_N FULL_COUNTER.COUNT_SUB_DFF10.Q 4.33e-19
C10568 sky130_fd_sc_hd__inv_1_6/Y FULL_COUNTER.COUNT_SUB_DFF1.Q 1.95e-20
C10569 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# V_GND 0.00228f
C10570 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.52e-19
C10571 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.00137f
C10572 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 5.13e-19
C10573 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 5.01e-19
C10574 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# V_LOW -0.313f
C10575 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# 5.29e-19
C10576 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00194f
C10577 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# sky130_fd_sc_hd__conb_1_28/HI -0.00581f
C10578 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_1_98/Y 0.00103f
C10579 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__inv_1_106/Y 0.0107f
C10580 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_57/Y 0.0277f
C10581 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_58/Y 0.00637f
C10582 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# -6.29e-19
C10583 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_557_413# -3.67e-20
C10584 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# -0.00126f
C10585 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# -7.77e-19
C10586 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# 0.00153f
C10587 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__nand3_1_2/B 3.24e-21
C10588 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 1.93e-21
C10589 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 2e-21
C10590 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 1.09e-20
C10591 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__conb_1_26/HI 0.00119f
C10592 sky130_fd_sc_hd__inv_1_5/Y V_GND 0.0841f
C10593 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -1.89e-19
C10594 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_31/a_473_413# 2.84e-32
C10595 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# -2.28e-19
C10596 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# V_LOW -7.25e-19
C10597 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# 0.00585f
C10598 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# V_GND -0.0466f
C10599 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF0.Q 5.66e-19
C10600 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# V_GND -0.0459f
C10601 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/Q_N 0.00391f
C10602 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# -0.00754f
C10603 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_557_413# -0.0012f
C10604 sky130_fd_sc_hd__inv_1_93/Y Reset 1.05e-19
C10605 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00136f
C10606 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__inv_1_9/Y 2.52e-19
C10607 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.3e-20
C10608 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# V_LOW 0.0254f
C10609 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.61e-19
C10610 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# V_LOW 4.8e-20
C10611 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__conb_1_26/HI 8.96e-21
C10612 sky130_fd_sc_hd__inv_1_46/A V_GND 0.12f
C10613 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.0194f
C10614 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 6.17e-19
C10615 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 8.11e-21
C10616 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# -1.76e-19
C10617 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 6.48e-20
C10618 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_97/Y 0.00132f
C10619 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# V_GND -0.0023f
C10620 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_119/Y 6.24e-21
C10621 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.47e-20
C10622 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.9e-19
C10623 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00412f
C10624 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__conb_1_39/HI -9.73e-19
C10625 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00471f
C10626 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.26e-20
C10627 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 8.26e-21
C10628 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# CLOCK_GEN.SR_Op.Q 7.52e-19
C10629 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# -2.65e-20
C10630 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 2.68e-21
C10631 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.92e-20
C10632 sky130_fd_sc_hd__inv_1_45/A V_GND 0.204f
C10633 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__inv_1_18/Y 0.0327f
C10634 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00544f
C10635 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_557_413# -3.67e-20
C10636 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# -0.00608f
C10637 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_381_47# 2.96e-20
C10638 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# V_LOW 1.26e-20
C10639 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# sky130_fd_sc_hd__inv_1_57/Y 0.00635f
C10640 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_18/HI 1.26e-19
C10641 sky130_fd_sc_hd__dfbbn_1_32/a_581_47# sky130_fd_sc_hd__inv_16_1/Y 0.00181f
C10642 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# -0.00458f
C10643 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_647_21# -0.00423f
C10644 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 5.07e-19
C10645 sky130_fd_sc_hd__dfbbn_1_42/a_581_47# V_GND 2.67e-19
C10646 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# V_LOW 1.79e-20
C10647 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00732f
C10648 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# V_GND 1.39e-19
C10649 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# V_LOW -2.68e-19
C10650 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__conb_1_35/HI 0.00121f
C10651 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# -0.05f
C10652 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 6.87e-20
C10653 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 9.38e-20
C10654 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 1.53e-19
C10655 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 5.62e-22
C10656 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__conb_1_40/HI 5.96e-19
C10657 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 4.85e-20
C10658 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__conb_1_30/HI 2.57e-20
C10659 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00739f
C10660 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF15.Q 8.34e-20
C10661 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.33e-20
C10662 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_16_1/Y 0.308f
C10663 FALLING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF7.Q 4.58e-19
C10664 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q -2.71e-20
C10665 sky130_fd_sc_hd__conb_1_34/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.197f
C10666 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# sky130_fd_sc_hd__nand3_1_0/Y 7.56e-19
C10667 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__inv_1_4/Y 1.3e-19
C10668 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# V_GND 1.64e-19
C10669 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# sky130_fd_sc_hd__conb_1_38/HI 0.00306f
C10670 sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# V_GND 1.11e-19
C10671 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 7.03e-19
C10672 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# 7.99e-20
C10673 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 9.52e-20
C10674 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_72/A 3.66e-19
C10675 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 0.0031f
C10676 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# sky130_fd_sc_hd__conb_1_28/HI 5.94e-19
C10677 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__conb_1_19/LO 0.0116f
C10678 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__conb_1_9/LO 6.16e-21
C10679 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_95/A 5.03e-20
C10680 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0156f
C10681 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# -1.66e-19
C10682 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.18e-20
C10683 Reset sky130_fd_sc_hd__inv_1_86/Y 0.00263f
C10684 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_70/A 0.0137f
C10685 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.00105f
C10686 sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__nand2_1_0/Y 0.00131f
C10687 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/Q_N -4.33e-20
C10688 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.19e-22
C10689 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# -0.0144f
C10690 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# -0.00431f
C10691 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__conb_1_17/HI -3.44e-19
C10692 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# -1.64e-19
C10693 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_8_5/a_27_47# 9.56e-20
C10694 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00108f
C10695 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# V_GND 2.85e-19
C10696 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 8.38e-21
C10697 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_64/A 0.052f
C10698 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 1.55e-19
C10699 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_2/HI 0.158f
C10700 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.84e-19
C10701 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# V_GND 2.39e-19
C10702 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# -5.42e-19
C10703 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_55/Y 0.024f
C10704 sky130_fd_sc_hd__nand3_1_0/a_109_47# sky130_fd_sc_hd__inv_1_66/Y 5.38e-19
C10705 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# V_LOW -0.32f
C10706 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 7e-20
C10707 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# V_LOW 0.0067f
C10708 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_32/HI 0.147f
C10709 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_557_413# -3.67e-20
C10710 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# -0.00946f
C10711 sky130_fd_sc_hd__nand3_1_0/a_109_47# V_GND -4.59e-19
C10712 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# 2.28e-19
C10713 sky130_fd_sc_hd__dfbbn_1_30/a_1112_329# sky130_fd_sc_hd__conb_1_40/HI 0.0015f
C10714 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 1.47e-21
C10715 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_647_21# 8.28e-20
C10716 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# V_GND -0.00397f
C10717 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0809f
C10718 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0436f
C10719 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__conb_1_16/HI 3.55e-20
C10720 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0163f
C10721 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.6e-19
C10722 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_39/HI -2.07e-19
C10723 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 5.72e-19
C10724 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# CLOCK_GEN.SR_Op.Q 2.03e-19
C10725 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 2.32e-20
C10726 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 1.45e-20
C10727 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 5.39e-20
C10728 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_100/Y 0.00455f
C10729 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.98e-21
C10730 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 1.21e-19
C10731 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# 1.86e-19
C10732 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 0.0395f
C10733 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__conb_1_18/HI 9.8e-19
C10734 sky130_fd_sc_hd__dfbbn_1_2/Q_N V_LOW -0.00509f
C10735 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_44/HI 3.11e-19
C10736 sky130_fd_sc_hd__inv_1_64/Y V_GND 0.0406f
C10737 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# V_GND -0.0408f
C10738 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# V_GND 0.00428f
C10739 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 9.88e-19
C10740 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_85/Y 0.00603f
C10741 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_17/LO 0.0134f
C10742 sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# sky130_fd_sc_hd__conb_1_32/HI 0.0049f
C10743 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# V_LOW 0.00676f
C10744 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.55e-19
C10745 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# sky130_fd_sc_hd__conb_1_35/HI 3.65e-19
C10746 sky130_fd_sc_hd__conb_1_36/HI V_LOW 0.147f
C10747 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__inv_1_112/Y 0.00192f
C10748 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0197f
C10749 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__conb_1_17/HI 3.69e-19
C10750 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_67/Y 1.63e-19
C10751 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF15.Q 0.029f
C10752 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.7e-20
C10753 sky130_fd_sc_hd__inv_1_72/Y V_GND 0.0573f
C10754 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00145f
C10755 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# sky130_fd_sc_hd__inv_1_5/Y 0.00315f
C10756 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.19e-20
C10757 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# -3.8e-20
C10758 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# -5.54e-21
C10759 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# -5.68e-32
C10760 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__inv_1_58/Y 0.0107f
C10761 FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_100/Y 0.00202f
C10762 sky130_fd_sc_hd__conb_1_47/HI sky130_fd_sc_hd__inv_1_108/Y 8.09e-20
C10763 sky130_fd_sc_hd__inv_1_56/Y sky130_fd_sc_hd__inv_16_0/Y 0.0115f
C10764 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__conb_1_36/LO 0.0102f
C10765 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 0.0127f
C10766 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# V_GND -0.00376f
C10767 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__nand2_1_2/A 1.91e-20
C10768 RISING_COUNTER.COUNT_SUB_DFF1.Q V_LOW 1.54f
C10769 sky130_fd_sc_hd__inv_1_119/Y V_SENSE 0.178f
C10770 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__conb_1_45/HI 5.11e-21
C10771 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__inv_1_7/Y 9.11e-20
C10772 sky130_fd_sc_hd__dfbbn_1_24/Q_N sky130_fd_sc_hd__conb_1_28/HI 2.64e-21
C10773 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 1.2e-20
C10774 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 2.58e-19
C10775 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 8.93e-20
C10776 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__conb_1_21/HI 4.51e-20
C10777 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_647_21# -0.00782f
C10778 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__nand3_1_2/Y 0.00158f
C10779 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_30/HI 0.00186f
C10780 sky130_fd_sc_hd__inv_1_61/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.103f
C10781 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# CLOCK_GEN.SR_Op.Q 2.8e-19
C10782 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 1.22e-19
C10783 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_26/HI 0.244f
C10784 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_16_1/Y 0.105f
C10785 sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.3e-19
C10786 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 0.0217f
C10787 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__conb_1_48/HI 5.85e-20
C10788 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# sky130_fd_sc_hd__inv_1_55/Y 7.87e-20
C10789 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0.0025f
C10790 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# -2.32e-19
C10791 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# -0.00147f
C10792 sky130_fd_sc_hd__conb_1_49/LO FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.01e-19
C10793 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# V_LOW -0.314f
C10794 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.2e-20
C10795 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 4.02e-19
C10796 sky130_fd_sc_hd__inv_1_42/Y V_GND 0.0758f
C10797 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__nand3_1_1/Y 0.0919f
C10798 sky130_fd_sc_hd__conb_1_39/HI Reset 3.11e-20
C10799 sky130_fd_sc_hd__conb_1_10/HI V_LOW 0.0411f
C10800 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_17/Y 0.365f
C10801 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 7.2e-21
C10802 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 2.29e-21
C10803 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 2.29e-21
C10804 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_581_47# 9.58e-20
C10805 sky130_fd_sc_hd__conb_1_42/LO FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.62e-20
C10806 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 1.2e-19
C10807 sky130_fd_sc_hd__dfbbn_1_0/Q_N V_GND -0.00693f
C10808 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00127f
C10809 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_24/LO 3.38e-21
C10810 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__conb_1_16/HI 8.93e-20
C10811 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0.00157f
C10812 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 1.53e-19
C10813 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 5.82e-19
C10814 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 1.68e-19
C10815 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0.00123f
C10816 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_13/LO 0.00122f
C10817 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__inv_1_102/Y 0.00565f
C10818 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.0432f
C10819 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# V_LOW 0.0128f
C10820 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.22e-19
C10821 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_4/HI 0.0372f
C10822 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__conb_1_2/HI 2.49e-19
C10823 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_1_18/Y 7.5e-19
C10824 RISING_COUNTER.COUNT_SUB_DFF5.Q V_LOW 5.32f
C10825 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 1.27e-19
C10826 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# V_GND -0.0105f
C10827 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 4.35e-19
C10828 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# 0.00145f
C10829 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# V_GND 1.58e-19
C10830 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# V_GND 0.0021f
C10831 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 0.00125f
C10832 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0199f
C10833 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_74/Y 0.0572f
C10834 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_381_47# 8.55e-21
C10835 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_75/Y 0.00542f
C10836 sky130_fd_sc_hd__dfbbn_1_41/a_581_47# sky130_fd_sc_hd__inv_1_112/Y 5.8e-19
C10837 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0352f
C10838 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__inv_1_107/Y 0.0491f
C10839 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# sky130_fd_sc_hd__nand3_1_2/Y 0.00136f
C10840 sky130_fd_sc_hd__nand2_1_3/Y V_LOW 0.00435f
C10841 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.62e-20
C10842 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.52e-20
C10843 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 6.09e-21
C10844 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_30/HI 0.186f
C10845 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__conb_1_0/HI 0.00498f
C10846 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# V_GND -0.0075f
C10847 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# sky130_fd_sc_hd__inv_1_103/Y 0.026f
C10848 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__conb_1_36/HI 0.00493f
C10849 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# -9.32e-20
C10850 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0246f
C10851 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__inv_1_61/Y 1.72e-20
C10852 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_6/LO 3.53e-19
C10853 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# V_GND -0.00493f
C10854 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# sky130_fd_sc_hd__conb_1_34/HI 1.57e-20
C10855 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.48e-19
C10856 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0727f
C10857 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 5.28e-19
C10858 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_38/HI 1e-18
C10859 FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_6/HI 0.177f
C10860 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# CLOCK_GEN.SR_Op.Q 8.11e-21
C10861 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__conb_1_24/HI 0.0106f
C10862 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.014f
C10863 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0055f
C10864 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 6.59e-20
C10865 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_581_47# -7.91e-19
C10866 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.34f
C10867 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__conb_1_2/HI 0.00451f
C10868 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# -1.69e-19
C10869 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__inv_1_102/Y 0.0686f
C10870 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.49e-21
C10871 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.734f
C10872 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_86/Y 0.00586f
C10873 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_67/Y 1.2e-19
C10874 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0.155f
C10875 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__conb_1_22/HI 0.0208f
C10876 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# sky130_fd_sc_hd__conb_1_49/LO 3.81e-20
C10877 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_8/HI 0.43f
C10878 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# 7.69e-20
C10879 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# sky130_fd_sc_hd__conb_1_48/HI 1.58e-19
C10880 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_16_2/Y 2.74e-19
C10881 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# 8.59e-20
C10882 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__conb_1_4/HI 3.65e-19
C10883 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_22/Y 6.43e-21
C10884 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 2.55e-19
C10885 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__inv_1_4/Y 0.00648f
C10886 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# -1.64e-19
C10887 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0389f
C10888 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# -7.17e-20
C10889 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00336f
C10890 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.56e-20
C10891 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_83/Y 2.05e-19
C10892 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# sky130_fd_sc_hd__conb_1_5/HI 0.00434f
C10893 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__conb_1_16/HI 9.8e-20
C10894 sky130_fd_sc_hd__conb_1_19/LO V_LOW 0.0653f
C10895 sky130_fd_sc_hd__dfbbn_1_25/Q_N RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0235f
C10896 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# V_LOW -0.00389f
C10897 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_891_329# 6.64e-20
C10898 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 8.67e-20
C10899 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_85/A 6.94e-19
C10900 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 2.96e-22
C10901 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/Q_N 4.16e-19
C10902 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 3.11e-19
C10903 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 2.96e-21
C10904 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.24e-19
C10905 sky130_fd_sc_hd__dfbbn_1_16/a_1340_413# sky130_fd_sc_hd__conb_1_4/HI 4.53e-19
C10906 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_1_100/Y 3.77e-20
C10907 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_27/LO 0.0143f
C10908 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_72/A 0.0429f
C10909 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 2.33e-19
C10910 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# V_GND 2.83e-19
C10911 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 1.28e-20
C10912 sky130_fd_sc_hd__inv_1_76/A V_LOW 1.43f
C10913 sky130_fd_sc_hd__dfbbn_1_41/Q_N V_GND -0.00762f
C10914 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# 4.48e-19
C10915 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 0.00978f
C10916 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# sky130_fd_sc_hd__inv_1_107/Y 0.0015f
C10917 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.0641f
C10918 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.00591f
C10919 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_10/HI 0.00171f
C10920 FALLING_COUNTER.COUNT_SUB_DFF12.Q V_LOW 2.54f
C10921 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.92e-19
C10922 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 0.0223f
C10923 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# V_GND 4.15e-19
C10924 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__conb_1_10/HI 4.97e-19
C10925 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# -9.52e-20
C10926 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__conb_1_44/LO 0.0143f
C10927 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__conb_1_0/HI 1.63e-20
C10928 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0.0012f
C10929 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# V_GND -0.0146f
C10930 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 5.07e-19
C10931 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.82e-20
C10932 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__conb_1_36/HI 0.0016f
C10933 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__inv_1_8/Y 0.0423f
C10934 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/Q_N -4.33e-20
C10935 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00674f
C10936 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.031f
C10937 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# sky130_fd_sc_hd__inv_1_61/Y 7.3e-20
C10938 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# sky130_fd_sc_hd__conb_1_11/HI 1.74e-19
C10939 sky130_fd_sc_hd__nand2_8_9/Y V_GND 0.0818f
C10940 sky130_fd_sc_hd__dfbbn_1_24/Q_N V_GND -0.00782f
C10941 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# sky130_fd_sc_hd__conb_1_34/HI -2.65e-20
C10942 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1_23/LO 7.32e-19
C10943 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0337f
C10944 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# sky130_fd_sc_hd__conb_1_42/HI 6.71e-19
C10945 sky130_fd_sc_hd__inv_1_13/Y V_LOW 0.0269f
C10946 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.0459f
C10947 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_10/Y 0.0246f
C10948 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# V_GND 0.00213f
C10949 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_581_47# 0.00187f
C10950 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.36e-19
C10951 FALLING_COUNTER.COUNT_SUB_DFF1.Q V_GND 1.38f
C10952 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_581_47# -7.91e-19
C10953 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_71/Y 0.00368f
C10954 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 3.67e-21
C10955 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 8e-21
C10956 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.22e-20
C10957 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00213f
C10958 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# V_GND 0.0369f
C10959 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.06e-21
C10960 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_20/Y 3.74e-20
C10961 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00184f
C10962 sky130_fd_sc_hd__inv_1_112/Y V_LOW 0.104f
C10963 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# V_GND -0.151f
C10964 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__inv_1_21/Y 0.0463f
C10965 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0277f
C10966 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# sky130_fd_sc_hd__conb_1_41/HI 3.12e-20
C10967 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__conb_1_34/HI 0.00466f
C10968 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 6.16e-21
C10969 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# sky130_fd_sc_hd__inv_1_20/Y 6.77e-20
C10970 sky130_fd_sc_hd__inv_1_64/A Reset 0.213f
C10971 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.77e-19
C10972 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.00287f
C10973 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# -0.00149f
C10974 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1112_329# 0.0026f
C10975 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.21e-20
C10976 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# sky130_fd_sc_hd__conb_1_5/HI 0.00207f
C10977 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.18e-20
C10978 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 7.69e-20
C10979 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF15.Q 0.311f
C10980 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_53/Y 2.37e-20
C10981 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.00109f
C10982 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_22/HI 0.00562f
C10983 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF19.Q 1.14f
C10984 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 3.31e-20
C10985 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 2.18e-19
C10986 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__conb_1_42/HI 0.00367f
C10987 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0323f
C10988 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# 3.61e-19
C10989 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 2.81e-19
C10990 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_22/Y 0.00147f
C10991 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00223f
C10992 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# V_GND -0.00149f
C10993 sky130_fd_sc_hd__inv_1_66/Y Reset 8.95e-21
C10994 sky130_fd_sc_hd__conb_1_25/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0545f
C10995 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# -0.0022f
C10996 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# -5.54e-21
C10997 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__inv_1_22/Y 2.3e-20
C10998 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 1.39e-19
C10999 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__inv_16_2/Y 5.11e-20
C11000 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.13e-19
C11001 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# V_LOW 1.38e-19
C11002 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.53e-19
C11003 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# V_LOW 0.0144f
C11004 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__conb_1_27/HI 0.00282f
C11005 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_791_47# 0.00126f
C11006 Reset V_GND 4.19f
C11007 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.29e-19
C11008 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 0.00488f
C11009 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__conb_1_10/HI -0.0088f
C11010 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_1_60/Y 0.00146f
C11011 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# V_LOW 0.00191f
C11012 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00136f
C11013 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# V_LOW -0.00121f
C11014 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_581_47# -2.6e-20
C11015 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_19/LO 5.58e-20
C11016 sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# sky130_fd_sc_hd__conb_1_36/HI 0.00138f
C11017 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_1_59/Y 0.0126f
C11018 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_47/HI -6.71e-19
C11019 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# 2.89e-19
C11020 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# 9e-21
C11021 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00116f
C11022 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 1.2e-19
C11023 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 0.00145f
C11024 sky130_fd_sc_hd__dfbbn_1_29/a_891_329# V_LOW 2.26e-20
C11025 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# V_GND 0.00207f
C11026 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# V_GND -0.04f
C11027 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# -5.54e-21
C11028 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# -0.00263f
C11029 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# V_LOW -3.29e-19
C11030 FALLING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF7.Q 5.26e-19
C11031 FULL_COUNTER.COUNT_SUB_DFF18.Q sky130_fd_sc_hd__inv_1_22/Y 0.35f
C11032 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# V_LOW 3.56e-20
C11033 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__nand3_1_1/Y 0.00384f
C11034 sky130_fd_sc_hd__inv_1_7/Y V_GND 0.181f
C11035 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# sky130_fd_sc_hd__inv_16_0/Y 8.67e-19
C11036 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# V_GND 0.00382f
C11037 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_1_58/Y 0.0149f
C11038 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 4.7e-19
C11039 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_6/Y 3.89e-20
C11040 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# V_GND -0.00479f
C11041 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_473_413# -3.86e-20
C11042 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_941_21# -1.61e-20
C11043 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 1.48e-19
C11044 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# V_LOW 0.00867f
C11045 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_41/HI 9.88e-20
C11046 FALLING_COUNTER.COUNT_SUB_DFF4.Q V_LOW 1.39f
C11047 sky130_fd_sc_hd__conb_1_18/LO V_LOW 0.0461f
C11048 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# V_GND 0.00653f
C11049 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 0.017f
C11050 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__conb_1_29/LO 1.88e-19
C11051 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__inv_16_2/Y 0.267f
C11052 sky130_fd_sc_hd__conb_1_11/LO V_GND -0.00325f
C11053 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 5.32e-19
C11054 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 6.55e-20
C11055 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 6.46e-20
C11056 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 0.00239f
C11057 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 0.00101f
C11058 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00119f
C11059 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 0.00621f
C11060 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# Reset 1.96e-19
C11061 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# V_GND 0.00345f
C11062 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_32/HI 5.28e-21
C11063 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_8_2/A 0.0218f
C11064 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# V_GND 3.34e-19
C11065 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# V_LOW 0.0106f
C11066 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_44/HI 0.0254f
C11067 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 9.17e-21
C11068 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# V_LOW 0.00712f
C11069 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# V_GND 2.23e-19
C11070 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# sky130_fd_sc_hd__inv_1_21/Y 3.1e-21
C11071 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# V_LOW 4.1e-19
C11072 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__nand2_8_0/a_27_47# 2.12e-19
C11073 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.18e-19
C11074 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.5e-19
C11075 sky130_fd_sc_hd__dfbbn_1_36/a_891_329# V_LOW -0.00121f
C11076 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.67e-20
C11077 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# V_GND -0.00188f
C11078 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_41/LO 1.21e-20
C11079 sky130_fd_sc_hd__dfbbn_1_48/Q_N RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0305f
C11080 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00767f
C11081 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 0.00105f
C11082 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# sky130_fd_sc_hd__inv_16_1/Y 1.37e-19
C11083 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__inv_1_16/Y 0.0219f
C11084 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__inv_1_101/Y 0.00231f
C11085 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_581_47# -2.6e-20
C11086 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF3.Q 5.11e-20
C11087 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 6.19e-19
C11088 sky130_fd_sc_hd__dfbbn_1_19/Q_N sky130_fd_sc_hd__conb_1_5/HI 3.16e-19
C11089 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_193_47# -0.228f
C11090 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.04e-19
C11091 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# Reset 0.0306f
C11092 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_62/Y 3.82e-21
C11093 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_32/HI 0.0243f
C11094 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 0.00942f
C11095 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 9.55e-19
C11096 Reset sky130_fd_sc_hd__nand3_1_1/Y 0.0669f
C11097 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# V_GND -0.0104f
C11098 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.299f
C11099 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__inv_1_60/Y 8.12e-20
C11100 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_21/Y 0.00213f
C11101 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# V_GND 0.00494f
C11102 FULL_COUNTER.COUNT_SUB_DFF6.Q V_GND 1.6f
C11103 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 9.36e-22
C11104 sky130_fd_sc_hd__inv_1_79/A V_LOW 0.162f
C11105 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# -2.3e-19
C11106 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# -0.0014f
C11107 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# V_GND 0.00119f
C11108 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# V_LOW 0.0111f
C11109 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 6.05e-19
C11110 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# V_GND -0.00475f
C11111 sky130_fd_sc_hd__inv_1_57/Y V_GND 0.0883f
C11112 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_25/LO 1.49e-19
C11113 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_5/HI 2.96e-20
C11114 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# -7.47e-20
C11115 sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 2.07e-19
C11116 sky130_fd_sc_hd__inv_1_17/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 9.87e-21
C11117 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0.00819f
C11118 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0302f
C11119 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0778f
C11120 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 6.07e-20
C11121 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# -5.54e-21
C11122 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# -0.00263f
C11123 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -2.6e-19
C11124 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_20/Y 9.69e-20
C11125 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 9.78e-19
C11126 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0.00738f
C11127 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 9.78e-19
C11128 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 1.03e-19
C11129 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 1.03e-19
C11130 sky130_fd_sc_hd__dfbbn_1_18/a_1363_47# sky130_fd_sc_hd__conb_1_9/HI -4.88e-19
C11131 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__conb_1_49/LO 2.09e-19
C11132 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_44/HI 0.272f
C11133 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_75/A 0.143f
C11134 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# V_LOW -0.00121f
C11135 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__conb_1_47/HI 0.00849f
C11136 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_16_1/Y 0.0999f
C11137 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# V_LOW 0.0107f
C11138 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_473_413# -5.33e-20
C11139 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# V_GND 0.00773f
C11140 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0177f
C11141 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__inv_1_12/Y 0.0337f
C11142 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_65/Y 0.0716f
C11143 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_13/HI 1.17e-21
C11144 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_12/Y 0.0298f
C11145 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__inv_1_12/Y 0.0119f
C11146 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# V_GND 2.64e-19
C11147 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_24/HI 2.55e-20
C11148 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# -9.32e-20
C11149 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 0.0332f
C11150 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.1e-21
C11151 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# -3.79e-20
C11152 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# -0.00336f
C11153 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 1.13e-19
C11154 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# V_GND 0.00186f
C11155 sky130_fd_sc_hd__inv_1_88/Y V_LOW 0.219f
C11156 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.73e-19
C11157 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__inv_1_58/Y 0.0238f
C11158 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# V_LOW 0.0444f
C11159 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0.431f
C11160 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_21/HI 1.37e-19
C11161 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_1_9/Y 0.0351f
C11162 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_38/HI 3.28e-19
C11163 sky130_fd_sc_hd__conb_1_28/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0148f
C11164 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# -2.57e-20
C11165 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 4.23e-19
C11166 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# -0.00729f
C11167 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_891_329# -1.42e-19
C11168 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_557_413# -0.0012f
C11169 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 2.63e-20
C11170 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 2.93e-20
C11171 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_32/HI 0.0316f
C11172 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__conb_1_26/LO 0.00206f
C11173 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# V_GND 0.00163f
C11174 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# V_LOW 0.00707f
C11175 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# V_GND -0.00401f
C11176 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_1_71/A 3.84e-19
C11177 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__conb_1_34/HI 1.03e-19
C11178 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 1.83e-22
C11179 sky130_fd_sc_hd__inv_1_54/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00128f
C11180 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_13/HI 1.26e-19
C11181 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.04e-20
C11182 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00404f
C11183 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.02e-21
C11184 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00106f
C11185 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# 2.09e-19
C11186 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_647_21# -6.43e-20
C11187 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_473_413# -0.00591f
C11188 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_36/LO 3.06e-21
C11189 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.08e-22
C11190 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.74e-20
C11191 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_557_413# 2.53e-19
C11192 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00552f
C11193 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.48e-20
C11194 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# V_GND -0.00465f
C11195 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF11.Q 0.129f
C11196 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.48e-20
C11197 sky130_fd_sc_hd__conb_1_37/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00544f
C11198 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.69e-19
C11199 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 2.26e-19
C11200 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# V_GND -0.0135f
C11201 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__conb_1_35/LO 8.81e-20
C11202 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 3.92e-19
C11203 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# Reset 0.0225f
C11204 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__conb_1_14/LO 7.06e-20
C11205 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 4.93e-19
C11206 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 2.86e-19
C11207 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00237f
C11208 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_85/Y 8.65e-20
C11209 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# V_GND -0.00732f
C11210 sky130_fd_sc_hd__conb_1_3/HI FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0739f
C11211 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_581_47# 5.8e-19
C11212 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 0.00739f
C11213 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# Reset 2.57e-20
C11214 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# 2.06e-20
C11215 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 3.72e-20
C11216 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.027f
C11217 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# 0.00228f
C11218 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.005f
C11219 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__conb_1_22/HI 0.00122f
C11220 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# V_GND 0.00203f
C11221 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_68/A 0.046f
C11222 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_70/A 0.131f
C11223 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/Q_N 0.00178f
C11224 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# -1.65e-19
C11225 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# -0.00591f
C11226 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_647_21# -6.43e-20
C11227 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_98/Y 6.46e-20
C11228 sky130_fd_sc_hd__conb_1_14/HI V_GND -0.0837f
C11229 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# V_GND 0.0015f
C11230 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_1_101/Y 8.59e-19
C11231 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# -2.37e-19
C11232 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_941_21# -3.07e-19
C11233 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 6.84e-21
C11234 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 0.00123f
C11235 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 1.68e-19
C11236 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0.00157f
C11237 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 1.53e-19
C11238 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 5.82e-19
C11239 sky130_fd_sc_hd__conb_1_42/HI sky130_fd_sc_hd__inv_1_103/Y 0.108f
C11240 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/Q_N -4.33e-20
C11241 sky130_fd_sc_hd__inv_1_68/A V_GND 0.17f
C11242 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -0.00139f
C11243 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# -2.3e-19
C11244 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.61e-19
C11245 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF0.Q 4.88e-19
C11246 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 7.66e-21
C11247 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# -9.32e-20
C11248 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# -5.54e-21
C11249 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# -0.00263f
C11250 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 1.33e-19
C11251 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.27e-20
C11252 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 1.07e-20
C11253 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 4.01e-20
C11254 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 4.01e-20
C11255 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00118f
C11256 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0113f
C11257 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 4.44e-20
C11258 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.0113f
C11259 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.00118f
C11260 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 4.44e-20
C11261 sky130_fd_sc_hd__inv_1_85/Y V_GND 0.0896f
C11262 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 7.65e-21
C11263 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00247f
C11264 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 5.6e-19
C11265 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 7.68e-20
C11266 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_11/LO 0.0141f
C11267 sky130_fd_sc_hd__conb_1_8/LO V_GND 0.00425f
C11268 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.00303f
C11269 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# V_LOW 1.79e-20
C11270 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_45/Y 0.00482f
C11271 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# -0.00255f
C11272 sky130_fd_sc_hd__inv_1_98/Y FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0261f
C11273 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/Q_N 0.00786f
C11274 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# V_GND 0.00593f
C11275 sky130_fd_sc_hd__dfbbn_1_12/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 4.52e-20
C11276 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__inv_16_1/Y 0.00148f
C11277 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__conb_1_22/HI 1.17e-21
C11278 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_40/HI 1.72e-20
C11279 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_23/Y 1.15e-19
C11280 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# sky130_fd_sc_hd__inv_1_12/Y 0.00913f
C11281 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# sky130_fd_sc_hd__inv_1_49/Y 0.00265f
C11282 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 4.45e-19
C11283 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/Q_N -4.24e-20
C11284 sky130_fd_sc_hd__dfbbn_1_11/Q_N V_LOW -0.0103f
C11285 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.3e-20
C11286 sky130_fd_sc_hd__inv_1_60/Y V_LOW 0.396f
C11287 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 2e-20
C11288 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_791_47# -5.42e-19
C11289 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 0.0451f
C11290 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# V_LOW 0.0043f
C11291 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__conb_1_39/HI 8.01e-21
C11292 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.59e-19
C11293 sky130_fd_sc_hd__dfbbn_1_12/Q_N V_GND 9.46e-19
C11294 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00199f
C11295 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__inv_1_9/Y 0.0458f
C11296 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_791_47# 0.00753f
C11297 sky130_fd_sc_hd__dfbbn_1_46/a_1340_413# V_LOW 2.94e-20
C11298 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 3.24e-20
C11299 sky130_fd_sc_hd__inv_1_28/Y V_GND 0.0843f
C11300 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_41/HI 0.0449f
C11301 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_45/A 0.0402f
C11302 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# -5.42e-19
C11303 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 4.53e-20
C11304 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__conb_1_32/HI 0.00725f
C11305 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__conb_1_26/LO 1.27e-19
C11306 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0307f
C11307 sky130_fd_sc_hd__inv_1_44/A V_LOW 0.0375f
C11308 sky130_fd_sc_hd__dfbbn_1_9/a_1363_47# V_GND -3.91e-19
C11309 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_70/A 1.6e-19
C11310 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_15/Y 2e-19
C11311 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 1.02e-19
C11312 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 1.02e-19
C11313 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# sky130_fd_sc_hd__conb_1_13/HI 1.61e-20
C11314 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_15/Y 0.205f
C11315 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 6.58e-20
C11316 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 3.44e-20
C11317 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0315f
C11318 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.31e-20
C11319 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 8.11e-21
C11320 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# V_GND 2.64e-19
C11321 sky130_fd_sc_hd__conb_1_35/LO Reset 0.014f
C11322 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# -0.0105f
C11323 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# -0.0193f
C11324 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# V_LOW 0.00556f
C11325 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# V_GND -0.00168f
C11326 sky130_fd_sc_hd__dfbbn_1_1/Q_N FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00103f
C11327 sky130_fd_sc_hd__inv_1_70/Y RISING_COUNTER.COUNT_SUB_DFF0.Q 4.4e-20
C11328 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 3.3e-20
C11329 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 1.59e-20
C11330 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# Reset 0.0108f
C11331 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 5.88e-21
C11332 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.83e-20
C11333 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.535f
C11334 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 8.63e-19
C11335 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 2.24e-20
C11336 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# V_GND -0.0131f
C11337 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_1159_47# 0.00225f
C11338 sky130_fd_sc_hd__inv_1_56/Y V_GND 0.0254f
C11339 sky130_fd_sc_hd__inv_1_68/A sky130_fd_sc_hd__nand3_1_1/Y 1.25e-19
C11340 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# -0.00548f
C11341 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_891_329# -0.00159f
C11342 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0278f
C11343 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00384f
C11344 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.00136f
C11345 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 4.17e-20
C11346 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_33/a_381_47# 8.67e-19
C11347 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0163f
C11348 sky130_fd_sc_hd__dfbbn_1_43/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.48e-19
C11349 sky130_fd_sc_hd__dfbbn_1_16/Q_N V_GND 0.00198f
C11350 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_31/LO 0.00154f
C11351 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# sky130_fd_sc_hd__inv_1_98/Y 3.34e-20
C11352 sky130_fd_sc_hd__dfbbn_1_14/Q_N V_GND -0.00245f
C11353 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# V_GND -0.00342f
C11354 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# sky130_fd_sc_hd__conb_1_51/HI 2.97e-19
C11355 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__conb_1_49/HI 0.0133f
C11356 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_891_329# 3.82e-21
C11357 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# -1.66e-19
C11358 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# -7.17e-20
C11359 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_80/A 3.96e-19
C11360 sky130_fd_sc_hd__inv_16_2/Y V_LOW 4.53f
C11361 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# V_LOW 0.00693f
C11362 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# 0.00629f
C11363 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 6.51e-19
C11364 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# -1.66e-19
C11365 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_43/A 9.63e-19
C11366 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_13/HI 0.0259f
C11367 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 1.36e-20
C11368 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 4.44e-20
C11369 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 2.44e-20
C11370 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 1.2e-19
C11371 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/Q_N -4.78e-20
C11372 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# -9.32e-20
C11373 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# V_LOW -0.00389f
C11374 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 2.96e-20
C11375 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00313f
C11376 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 2.96e-20
C11377 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_2_0/Y 3.24e-20
C11378 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_381_47# -0.00889f
C11379 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# -8.96e-20
C11380 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# -6.23e-21
C11381 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_791_47# 3.45e-20
C11382 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 9.22e-20
C11383 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_1_20/Y 0.00105f
C11384 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__inv_1_67/Y 1.22e-20
C11385 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_75/A 1.16e-20
C11386 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_17/HI 1.86e-20
C11387 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# V_LOW 0.0171f
C11388 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# CLOCK_GEN.SR_Op.Q 5.97e-21
C11389 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__inv_1_13/Y 1.5e-20
C11390 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__inv_1_8/Y 1.72e-20
C11391 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# V_LOW 0.00743f
C11392 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# V_GND 0.00256f
C11393 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 2.49e-19
C11394 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_20/HI 0.43f
C11395 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_45/LO 0.0702f
C11396 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_1_12/Y 0.00156f
C11397 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_891_329# 6.89e-19
C11398 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 0.00111f
C11399 FALLING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_108/Y 0.0111f
C11400 sky130_fd_sc_hd__inv_1_119/Y sky130_fd_sc_hd__inv_2_0/A 0.185f
C11401 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# V_LOW -0.00325f
C11402 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.23e-19
C11403 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__conb_1_39/HI 7.89e-21
C11404 sky130_fd_sc_hd__dfbbn_1_25/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0109f
C11405 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_57/Y 7.34e-21
C11406 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# V_GND 5.05e-19
C11407 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_41/HI 0.0409f
C11408 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__inv_1_90/Y 0.00547f
C11409 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 6.84e-22
C11410 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 5.82e-21
C11411 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0.00453f
C11412 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00553f
C11413 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 0.00305f
C11414 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# V_GND 0.00151f
C11415 sky130_fd_sc_hd__inv_1_102/Y sky130_fd_sc_hd__inv_16_1/Y 0.537f
C11416 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 0.00388f
C11417 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_18/LO 8.9e-21
C11418 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# V_GND 4.54e-19
C11419 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__inv_1_15/Y 0.00507f
C11420 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0135f
C11421 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.00453f
C11422 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_1/Y 3.47e-19
C11423 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 0.00559f
C11424 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_1_16/Y 2.15e-19
C11425 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__inv_1_103/Y 0.00379f
C11426 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 4.06e-21
C11427 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_16_1/Y 4.82e-22
C11428 RISING_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 6.82e-19
C11429 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 6.71e-19
C11430 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 3.27e-20
C11431 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_91/Y 0.0331f
C11432 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 6.95e-20
C11433 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/Q_N 4.77e-20
C11434 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# -0.0144f
C11435 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_647_21# -0.0106f
C11436 sky130_fd_sc_hd__conb_1_30/HI V_GND -0.12f
C11437 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__inv_1_61/Y 0.00153f
C11438 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0.00298f
C11439 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 1.77f
C11440 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 2.61e-19
C11441 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.06e-21
C11442 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 5.88e-19
C11443 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 0.00863f
C11444 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 7.67e-19
C11445 sky130_fd_sc_hd__dfbbn_1_3/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.1e-19
C11446 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 5.77e-20
C11447 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 9.7e-21
C11448 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__conb_1_35/HI 0.0368f
C11449 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# Reset 0.00135f
C11450 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 7.3e-20
C11451 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__conb_1_45/HI 4.1e-19
C11452 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 6.07e-19
C11453 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# -3.46e-20
C11454 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 2.29e-19
C11455 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 0.00185f
C11456 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.72e-20
C11457 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_80/A 6.08e-20
C11458 sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__inv_1_93/A 4.06e-21
C11459 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 3.78e-19
C11460 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 7.97e-19
C11461 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.3e-21
C11462 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0272f
C11463 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__inv_1_23/Y 0.0107f
C11464 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 9.69e-22
C11465 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# V_GND -0.00509f
C11466 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0406f
C11467 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.99e-20
C11468 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 1.69e-19
C11469 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0.00131f
C11470 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 1.78e-19
C11471 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 1.32e-19
C11472 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 6.03e-19
C11473 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.271f
C11474 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0727f
C11475 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# 2.3e-19
C11476 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0324f
C11477 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 7.48e-19
C11478 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 3.24e-19
C11479 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 3.55e-20
C11480 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00225f
C11481 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 1.91e-19
C11482 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 9.29e-21
C11483 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.1e-19
C11484 FALLING_COUNTER.COUNT_SUB_DFF3.Q V_LOW 1.19f
C11485 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/Q_N -4.24e-20
C11486 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__conb_1_46/HI -2.59e-19
C11487 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__conb_1_2/HI 8.1e-20
C11488 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_17/HI 1.72e-20
C11489 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/Q_N 5.85e-22
C11490 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0894f
C11491 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# sky130_fd_sc_hd__inv_1_103/Y 0.00269f
C11492 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__inv_1_20/Y 4.07e-20
C11493 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__conb_1_35/LO 4.54e-20
C11494 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# V_LOW 1.79e-20
C11495 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__conb_1_47/HI 3.89e-19
C11496 sky130_fd_sc_hd__fill_4_84/VPB V_LOW 0.797f
C11497 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__inv_1_15/Y 5.37e-20
C11498 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# V_LOW -2.78e-35
C11499 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# V_GND 0.00214f
C11500 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 6.25e-21
C11501 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 1.49e-20
C11502 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 3.07e-19
C11503 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 5.15e-19
C11504 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 5.56e-19
C11505 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 4.79e-19
C11506 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 3.21e-20
C11507 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 3.2e-20
C11508 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.14e-19
C11509 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_557_413# 0.00136f
C11510 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.0278f
C11511 sky130_fd_sc_hd__conb_1_29/HI RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0136f
C11512 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__conb_1_39/HI 6.57e-20
C11513 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# V_LOW 0.0166f
C11514 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 5.44e-20
C11515 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_16_0/Y 0.898f
C11516 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 0.352f
C11517 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 5.36e-19
C11518 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 3.8e-21
C11519 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# V_LOW 0.0122f
C11520 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 5.22e-19
C11521 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_1_112/Y 0.0098f
C11522 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0891f
C11523 sky130_fd_sc_hd__inv_1_96/A V_LOW 0.355f
C11524 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.0595f
C11525 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# V_LOW 0.00263f
C11526 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 3.87e-20
C11527 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__inv_1_13/Y 2.78e-20
C11528 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 6.81e-19
C11529 sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# V_GND 1.64e-19
C11530 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 1.02f
C11531 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.00249f
C11532 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_891_329# -3.85e-20
C11533 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# -4.1e-19
C11534 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0929f
C11535 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.9e-20
C11536 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_54/Y 0.0011f
C11537 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__conb_1_6/HI 8.48e-20
C11538 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# 2.88e-19
C11539 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 2.88e-19
C11540 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00776f
C11541 sky130_fd_sc_hd__dfbbn_1_10/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00721f
C11542 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# sky130_fd_sc_hd__inv_1_16/Y 2.14e-20
C11543 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 4.03e-19
C11544 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 7.16e-19
C11545 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 5.68e-20
C11546 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 7.16e-19
C11547 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 4.03e-19
C11548 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 5.68e-20
C11549 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# V_LOW 0.0332f
C11550 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_11/Y 1.19e-19
C11551 sky130_fd_sc_hd__conb_1_32/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00395f
C11552 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# V_GND -0.00434f
C11553 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# V_GND 0.00131f
C11554 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# sky130_fd_sc_hd__conb_1_22/HI 3.63e-20
C11555 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_193_47# -0.0127f
C11556 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_36/LO 0.00216f
C11557 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0.557f
C11558 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# V_GND 0.00155f
C11559 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.102f
C11560 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# V_GND 0.00641f
C11561 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_40/a_381_47# 0.0124f
C11562 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.00209f
C11563 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# V_GND 0.00348f
C11564 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 0.00243f
C11565 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# 3.1e-19
C11566 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# sky130_fd_sc_hd__conb_1_35/HI 9.52e-19
C11567 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF13.Q 0.146f
C11568 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_1_23/Y 1.18e-19
C11569 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_96/Y 0.00141f
C11570 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 1.65e-19
C11571 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF14.Q 4.43e-21
C11572 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# sky130_fd_sc_hd__conb_1_45/HI 0.00115f
C11573 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# sky130_fd_sc_hd__inv_16_1/Y 1.14e-19
C11574 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.31e-20
C11575 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.22e-20
C11576 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0194f
C11577 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.94e-21
C11578 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__conb_1_49/HI 0.00162f
C11579 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__conb_1_0/HI 6.41e-19
C11580 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# V_GND 0.00263f
C11581 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# V_GND 0.0177f
C11582 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 1.55e-19
C11583 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 1e-18
C11584 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00473f
C11585 sky130_fd_sc_hd__dfbbn_1_49/Q_N V_GND -0.0074f
C11586 sky130_fd_sc_hd__conb_1_25/LO V_LOW 0.0818f
C11587 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# 1.34e-20
C11588 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0.00106f
C11589 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0249f
C11590 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 0.0106f
C11591 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__conb_1_9/HI 0.0229f
C11592 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__inv_1_11/Y 3.81e-19
C11593 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 2.9e-19
C11594 sky130_fd_sc_hd__conb_1_32/LO V_LOW 0.0809f
C11595 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00173f
C11596 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_16_1/Y 4.85e-21
C11597 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# V_LOW 0.043f
C11598 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_102/Y 3.54e-19
C11599 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# 7.63e-20
C11600 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# 5.26e-21
C11601 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0475f
C11602 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0576f
C11603 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_791_47# 8.23e-19
C11604 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 1.31e-19
C11605 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0434f
C11606 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 5.12e-21
C11607 sky130_fd_sc_hd__dfbbn_1_1/a_1363_47# sky130_fd_sc_hd__conb_1_2/HI -2.65e-20
C11608 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# -3.48e-20
C11609 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_891_329# -2.2e-20
C11610 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0426f
C11611 FALLING_COUNTER.COUNT_SUB_DFF12.Q FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0196f
C11612 sky130_fd_sc_hd__conb_1_43/LO V_LOW 0.103f
C11613 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/Q_N -9.56e-20
C11614 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 1.28e-19
C11615 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.373f
C11616 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__inv_1_20/Y 1.72e-20
C11617 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_86/Y 0.176f
C11618 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_56/Y 0.159f
C11619 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 9.49e-21
C11620 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# sky130_fd_sc_hd__conb_1_47/HI 1.14e-19
C11621 sky130_fd_sc_hd__dfbbn_1_3/Q_N V_LOW -0.00141f
C11622 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__conb_1_24/HI 9.87e-21
C11623 sky130_fd_sc_hd__dfbbn_1_17/Q_N V_GND 0.00258f
C11624 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# -8.61e-20
C11625 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# V_GND -0.00322f
C11626 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__inv_1_11/Y 0.0454f
C11627 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.84e-20
C11628 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 7.55e-20
C11629 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_99/Y 3.19e-21
C11630 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.79e-20
C11631 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__conb_1_39/HI 2.25e-19
C11632 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# V_LOW 2.94e-20
C11633 sky130_fd_sc_hd__dfbbn_1_26/a_891_329# V_LOW -0.00121f
C11634 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 8.26e-21
C11635 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_1112_329# 1.65e-19
C11636 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 7.2e-20
C11637 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__inv_1_17/Y 9.9e-19
C11638 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_18/Y 0.182f
C11639 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 8.58e-19
C11640 RISING_COUNTER.COUNT_SUB_DFF15.Q V_GND 0.899f
C11641 sky130_fd_sc_hd__conb_1_29/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.76e-20
C11642 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# V_LOW 1.79e-20
C11643 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 7.31e-21
C11644 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 2.11e-20
C11645 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF9.Q 1.04e-19
C11646 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.16e-20
C11647 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# V_LOW 2.26e-20
C11648 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_557_413# -0.0012f
C11649 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# -0.019f
C11650 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_1_100/Y 1.53e-20
C11651 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00178f
C11652 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# sky130_fd_sc_hd__inv_16_1/Y 0.00159f
C11653 sky130_fd_sc_hd__dfbbn_1_45/a_1340_413# V_LOW -6.55e-19
C11654 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 5.12e-19
C11655 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# 2.66e-19
C11656 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# -0.00385f
C11657 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.00391f
C11658 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__inv_1_54/Y 0.00141f
C11659 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_72/A 4.54e-19
C11660 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 3.87e-19
C11661 sky130_fd_sc_hd__dfbbn_1_21/Q_N RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0295f
C11662 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_42/HI 0.555f
C11663 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0.00135f
C11664 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 0.00135f
C11665 sky130_fd_sc_hd__dfbbn_1_18/a_1340_413# V_LOW 2.94e-20
C11666 V_GND V_HIGH 31.4f
C11667 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_17/Y 0.0163f
C11668 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# V_GND -0.0015f
C11669 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# V_GND -0.0046f
C11670 sky130_fd_sc_hd__dfbbn_1_44/a_557_413# V_LOW 3.56e-20
C11671 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_105/Y 0.0511f
C11672 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_67/Y 0.00358f
C11673 sky130_fd_sc_hd__dfbbn_1_15/a_1363_47# V_GND 1.46e-19
C11674 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_1_99/Y 0.0125f
C11675 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 2.88e-19
C11676 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# V_GND 0.00177f
C11677 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0104f
C11678 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__conb_1_25/HI 6.18e-19
C11679 sky130_fd_sc_hd__inv_1_9/Y V_LOW 0.402f
C11680 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 8.84e-19
C11681 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# V_GND 6.11e-19
C11682 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# V_LOW 0.0103f
C11683 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 0.00222f
C11684 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# V_GND 0.0202f
C11685 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# -0.00144f
C11686 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_80/A 0.0701f
C11687 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__inv_1_23/Y 2.42e-19
C11688 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_19/Q_N 3.15e-20
C11689 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 6.1e-19
C11690 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_83/Y 0.0046f
C11691 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 1.51f
C11692 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0932f
C11693 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_381_47# -0.00144f
C11694 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.12e-20
C11695 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_891_329# 4.06e-19
C11696 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# sky130_fd_sc_hd__conb_1_49/HI 4.31e-19
C11697 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# sky130_fd_sc_hd__conb_1_0/HI 0.0017f
C11698 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_78/A 3.79e-20
C11699 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# V_GND -0.00146f
C11700 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_2_0/Y 8.5e-19
C11701 sky130_fd_sc_hd__dfbbn_1_42/a_891_329# sky130_fd_sc_hd__inv_1_59/Y 5.46e-20
C11702 FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__nand3_1_2/B 4.06e-21
C11703 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# V_GND 1.48e-19
C11704 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 3.27e-20
C11705 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 2.25e-20
C11706 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# Reset 0.0221f
C11707 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.84e-20
C11708 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00261f
C11709 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0161f
C11710 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__inv_16_2/Y 0.0111f
C11711 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/Q_N 2.66e-19
C11712 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 0.00146f
C11713 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# 7.89e-19
C11714 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_50/A 0.0462f
C11715 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.054f
C11716 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# -0.00478f
C11717 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_16_0/Y 0.224f
C11718 sky130_fd_sc_hd__conb_1_6/HI V_GND 0.109f
C11719 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# V_GND 0.00166f
C11720 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# V_LOW -6.55e-19
C11721 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.00824f
C11722 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_1_19/Y 6.84e-19
C11723 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# -1.89e-19
C11724 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# -2.32e-19
C11725 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_791_47# 7.89e-19
C11726 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.218f
C11727 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0549f
C11728 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 3.14e-21
C11729 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 3.14e-21
C11730 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.3e-19
C11731 sky130_fd_sc_hd__dfbbn_1_33/Q_N FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.91e-19
C11732 sky130_fd_sc_hd__nand3_1_2/B V_LOW 0.136f
C11733 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_10/Y 1.21e-19
C11734 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0191f
C11735 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 4.78e-19
C11736 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 4.78e-19
C11737 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# -0.00142f
C11738 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.0293f
C11739 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# -5.33e-20
C11740 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_557_413# -3.67e-20
C11741 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__inv_1_21/Y 2.95e-19
C11742 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 1.32e-20
C11743 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 0.00523f
C11744 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_94/A 5.11e-19
C11745 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__conb_1_2/HI 0.00191f
C11746 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.84e-20
C11747 sky130_fd_sc_hd__inv_1_102/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00446f
C11748 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_47/HI 1.43e-20
C11749 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_54/Y 7.14e-20
C11750 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_16/HI 0.00553f
C11751 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__conb_1_35/HI 1.74e-20
C11752 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_581_47# -7.91e-19
C11753 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# V_GND 6.07e-19
C11754 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# sky130_fd_sc_hd__inv_1_11/Y 0.00156f
C11755 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF11.Q 0.156f
C11756 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_70/A 0.0527f
C11757 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_54/Y 0.00177f
C11758 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# -0.00379f
C11759 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 7.62e-20
C11760 sky130_fd_sc_hd__inv_1_49/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.379f
C11761 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# sky130_fd_sc_hd__inv_1_17/Y 1.04e-19
C11762 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_37/LO 0.012f
C11763 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# -0.00519f
C11764 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0098f
C11765 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# V_LOW -4.03e-19
C11766 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.102f
C11767 sky130_fd_sc_hd__inv_1_102/Y V_LOW 0.359f
C11768 sky130_fd_sc_hd__inv_1_12/Y sky130_fd_sc_hd__conb_1_6/HI 0.0193f
C11769 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# -5.42e-19
C11770 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 9.3e-21
C11771 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# V_LOW -0.00121f
C11772 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 4.62e-19
C11773 FULL_COUNTER.COUNT_SUB_DFF13.Q V_LOW 1.87f
C11774 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.0601f
C11775 sky130_fd_sc_hd__inv_1_49/Y V_LOW 0.363f
C11776 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.38e-21
C11777 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_59/Y 2.21e-20
C11778 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.00497f
C11779 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_17/HI 0.0107f
C11780 sky130_fd_sc_hd__dfbbn_1_31/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 8.26e-19
C11781 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_791_47# 3.56e-20
C11782 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 3.56e-20
C11783 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__conb_1_25/HI 0.0231f
C11784 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0057f
C11785 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0205f
C11786 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 7.96e-21
C11787 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 0.0107f
C11788 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# V_GND 2.67e-20
C11789 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 9.02e-19
C11790 FULL_COUNTER.COUNT_SUB_DFF17.Q V_GND 2.85f
C11791 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__conb_1_21/HI 4.38e-19
C11792 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_1_11/Y 0.0103f
C11793 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_97/A 0.00449f
C11794 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.0024f
C11795 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# V_LOW 0.00914f
C11796 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# -7.77e-19
C11797 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# -0.00115f
C11798 sky130_fd_sc_hd__conb_1_29/LO sky130_fd_sc_hd__inv_1_59/Y 0.0305f
C11799 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00372f
C11800 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# -1.44e-20
C11801 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# V_LOW 1.79e-20
C11802 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# V_GND 0.0016f
C11803 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 0.00334f
C11804 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 9.72e-19
C11805 sky130_fd_sc_hd__inv_1_33/Y V_SENSE 0.147f
C11806 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00395f
C11807 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 1.42e-20
C11808 sky130_fd_sc_hd__dfbbn_1_2/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00102f
C11809 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# -0.00141f
C11810 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 3.13e-20
C11811 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# -2.02e-19
C11812 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# -5.54e-21
C11813 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.00896f
C11814 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 1.33e-19
C11815 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0676f
C11816 sky130_fd_sc_hd__conb_1_50/LO RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0495f
C11817 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_19/Y 0.189f
C11818 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_473_413# 6.75e-20
C11819 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# 2.6e-20
C11820 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# Reset 0.0171f
C11821 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 8.94e-20
C11822 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_26/HI 0.126f
C11823 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.34e-20
C11824 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 6.95e-20
C11825 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__inv_16_0/Y 0.0222f
C11826 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 0.00209f
C11827 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0472f
C11828 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# V_GND 0.0118f
C11829 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00151f
C11830 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_581_47# -7.91e-19
C11831 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# V_GND 1.48e-19
C11832 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# -1.64e-19
C11833 sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 0.00218f
C11834 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 7.3e-22
C11835 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__inv_1_57/Y 3.49e-19
C11836 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__conb_1_20/HI -0.00229f
C11837 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0365f
C11838 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 6.64e-20
C11839 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 6.64e-20
C11840 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_93/A 0.0261f
C11841 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0192f
C11842 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_24/LO 8.84e-20
C11843 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 5.57e-22
C11844 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_381_47# -0.00527f
C11845 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# -6.23e-21
C11846 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# CLOCK_GEN.SR_Op.Q 5.71e-19
C11847 sky130_fd_sc_hd__conb_1_34/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0497f
C11848 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 4.43e-21
C11849 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# sky130_fd_sc_hd__conb_1_2/HI 3.8e-19
C11850 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__inv_1_59/Y 1.4e-21
C11851 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# -4.66e-20
C11852 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# sky130_fd_sc_hd__dfbbn_1_3/a_381_47# -3.79e-20
C11853 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 8.66e-21
C11854 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 4.44e-20
C11855 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 6.4e-19
C11856 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 1.08e-19
C11857 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_581_47# -7.91e-19
C11858 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.29e-19
C11859 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_86/Y 8.33e-20
C11860 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__inv_1_55/Y 2.85e-20
C11861 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# V_LOW 0.033f
C11862 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0242f
C11863 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_581_47# -7.91e-19
C11864 sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00222f
C11865 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0238f
C11866 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 0.0027f
C11867 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 8.19e-21
C11868 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_1/LO 9.27e-19
C11869 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# sky130_fd_sc_hd__inv_1_11/Y 1.44e-19
C11870 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_31/HI 6.04e-19
C11871 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 7.07e-19
C11872 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.87e-20
C11873 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.59e-20
C11874 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__inv_1_119/Y 5.29e-20
C11875 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 4.63e-23
C11876 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 8.6e-23
C11877 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.85e-21
C11878 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# sky130_fd_sc_hd__inv_1_90/Y 3.75e-21
C11879 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00107f
C11880 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# sky130_fd_sc_hd__inv_1_9/Y 5.62e-19
C11881 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# V_GND -0.00199f
C11882 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00263f
C11883 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.91e-19
C11884 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# V_GND 0.00367f
C11885 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__conb_1_21/HI 0.00117f
C11886 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__inv_1_11/Y 1.53e-19
C11887 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0301f
C11888 sky130_fd_sc_hd__dfbbn_1_17/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 1.12e-19
C11889 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# V_LOW 1.07e-19
C11890 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# -1.66e-19
C11891 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 3.41e-20
C11892 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_45/HI 0.0224f
C11893 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 7.89e-19
C11894 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 0.00115f
C11895 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_1340_413# 1.1e-19
C11896 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__inv_1_106/Y 3.19e-19
C11897 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 3.76e-21
C11898 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_71/Y 0.27f
C11899 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 4.76e-19
C11900 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00198f
C11901 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__inv_16_2/Y 2.53e-20
C11902 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 0.00821f
C11903 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 1.04f
C11904 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 3.18e-20
C11905 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 4.5e-19
C11906 RISING_COUNTER.COUNT_SUB_DFF8.Q RISING_COUNTER.COUNT_SUB_DFF5.Q 2.34e-19
C11907 sky130_fd_sc_hd__dfbbn_1_46/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.38e-19
C11908 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.28e-19
C11909 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# -9.32e-20
C11910 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.00616f
C11911 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 3e-21
C11912 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.74e-21
C11913 sky130_fd_sc_hd__inv_1_74/Y V_LOW 0.222f
C11914 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0369f
C11915 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 8.28e-20
C11916 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 8.99e-20
C11917 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__conb_1_5/HI 8.63e-20
C11918 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0848f
C11919 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# V_GND 0.00488f
C11920 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__conb_1_20/HI -1.64e-19
C11921 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 6.17e-19
C11922 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 6.79e-21
C11923 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 2.2e-19
C11924 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.00283f
C11925 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF13.Q 2.53e-20
C11926 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 0.429f
C11927 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 8.74e-21
C11928 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 8.48e-21
C11929 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.00571f
C11930 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_44/HI 1.62e-19
C11931 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 3.42e-20
C11932 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__conb_1_41/LO 7.01e-20
C11933 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_16/HI 1.01e-20
C11934 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_1363_47# 6.52e-20
C11935 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 7.67e-19
C11936 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 8.83e-19
C11937 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 5.03e-19
C11938 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.04e-20
C11939 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# 1.67e-19
C11940 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__conb_1_23/HI -0.0185f
C11941 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.42e-20
C11942 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# sky130_fd_sc_hd__inv_1_55/Y 7.69e-22
C11943 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_54/Y 0.099f
C11944 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 0.00115f
C11945 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 1.27e-19
C11946 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.34e-20
C11947 sky130_fd_sc_hd__dfbbn_1_39/a_1340_413# V_LOW -6.55e-19
C11948 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__inv_1_53/Y 8.7e-20
C11949 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 2.3e-22
C11950 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__nand2_8_2/A 5.38e-20
C11951 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 0.00131f
C11952 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_25/HI 0.0892f
C11953 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 1.24e-20
C11954 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.00377f
C11955 FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_15/Y 3.17e-20
C11956 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0959f
C11957 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.036f
C11958 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_581_47# 3.11e-20
C11959 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.5e-19
C11960 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_101/Y -0.00108f
C11961 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00135f
C11962 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# 1.52e-19
C11963 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00153f
C11964 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.84e-22
C11965 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.09e-19
C11966 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 6.89e-21
C11967 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_20/Y 0.0268f
C11968 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.27e-19
C11969 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# V_LOW -5.87e-19
C11970 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# CLOCK_GEN.SR_Op.Q 0.0353f
C11971 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__conb_1_12/HI 4.89e-19
C11972 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 4.88e-20
C11973 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 3.48e-19
C11974 sky130_fd_sc_hd__dfbbn_1_11/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00172f
C11975 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.12e-19
C11976 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_76/A 5.5e-20
C11977 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# V_GND 6.67e-19
C11978 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_1_105/Y 0.0081f
C11979 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_75/A 0.00737f
C11980 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_53/Y 0.114f
C11981 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__inv_1_54/Y 0.0666f
C11982 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_1_11/Y 0.00317f
C11983 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 2.27e-19
C11984 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 7.9e-19
C11985 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 1.62e-19
C11986 FALLING_COUNTER.COUNT_SUB_DFF2.Q FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.08f
C11987 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__conb_1_31/HI 3.94e-21
C11988 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_76/A 9.92e-20
C11989 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_6/LO 3.75e-21
C11990 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0.00122f
C11991 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__conb_1_26/HI 1.22e-20
C11992 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 1.69e-20
C11993 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# sky130_fd_sc_hd__conb_1_37/HI -2.65e-20
C11994 sky130_fd_sc_hd__conb_1_43/HI FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0235f
C11995 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.0044f
C11996 FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_101/Y 0.124f
C11997 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 9.55e-19
C11998 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.82e-19
C11999 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0359f
C12000 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1363_47# 2.29e-19
C12001 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__inv_1_18/Y 5.95e-19
C12002 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.00237f
C12003 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 2.45e-19
C12004 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 1.19e-20
C12005 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_6/HI -0.00122f
C12006 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 4.7e-21
C12007 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# V_GND 3.96e-19
C12008 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/Q_N -4.33e-20
C12009 sky130_fd_sc_hd__inv_1_89/Y V_GND 0.0349f
C12010 sky130_fd_sc_hd__dfbbn_1_5/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00224f
C12011 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__conb_1_0/HI 0.00301f
C12012 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0304f
C12013 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 2.1e-19
C12014 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0048f
C12015 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__conb_1_5/HI 1.82e-20
C12016 sky130_fd_sc_hd__inv_1_52/Y V_LOW 0.2f
C12017 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_94/A 0.0302f
C12018 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 0.00575f
C12019 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_11/HI 0.189f
C12020 sky130_fd_sc_hd__nand3_1_2/Y V_GND 0.194f
C12021 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.387f
C12022 FULL_COUNTER.COUNT_SUB_DFF9.Q FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0825f
C12023 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 3.41e-19
C12024 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__conb_1_21/HI 0.0142f
C12025 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# sky130_fd_sc_hd__conb_1_28/HI 3.38e-21
C12026 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__inv_1_99/Y 4.77e-21
C12027 sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 0.00101f
C12028 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.00162f
C12029 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 6.47e-19
C12030 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.0037f
C12031 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 1.08e-20
C12032 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 2.82e-20
C12033 FULL_COUNTER.COUNT_SUB_DFF15.Q CLOCK_GEN.SR_Op.Q 0.3f
C12034 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# -0.00782f
C12035 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 9.63e-22
C12036 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# -1.38e-19
C12037 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# -5.54e-21
C12038 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# sky130_fd_sc_hd__conb_1_44/HI 1.85e-19
C12039 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0147f
C12040 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_1_98/Y 0.0596f
C12041 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.61e-20
C12042 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__conb_1_18/HI 8.14e-20
C12043 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__inv_16_2/Y 0.91f
C12044 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# sky130_fd_sc_hd__inv_1_58/Y 2.45e-20
C12045 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.23e-20
C12046 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_80/A 0.0388f
C12047 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0012f
C12048 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__conb_1_28/LO 8.84e-20
C12049 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 0.03f
C12050 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__conb_1_1/LO 8.84e-20
C12051 sky130_fd_sc_hd__conb_1_49/HI V_GND 0.106f
C12052 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.75e-19
C12053 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__conb_1_2/HI 1.66e-20
C12054 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 2.87e-20
C12055 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_21/Y 1.7e-19
C12056 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 7.23e-21
C12057 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 8.6e-21
C12058 sky130_fd_sc_hd__conb_1_51/LO sky130_fd_sc_hd__conb_1_38/HI 1.73e-20
C12059 sky130_fd_sc_hd__inv_1_59/Y V_LOW 0.199f
C12060 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0.0682f
C12061 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 1.38e-20
C12062 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__nand3_1_2/B 8.66e-20
C12063 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__conb_1_30/HI -0.00143f
C12064 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# -6.23e-21
C12065 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# -4.5e-20
C12066 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__inv_1_106/Y 0.0155f
C12067 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# V_LOW -2.78e-35
C12068 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 9.24e-21
C12069 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0.0388f
C12070 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.85e-21
C12071 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 5.45e-22
C12072 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 2.89e-20
C12073 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 3.12e-21
C12074 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_22/HI 0.0256f
C12075 sky130_fd_sc_hd__conb_1_4/LO sky130_fd_sc_hd__inv_16_2/Y 8.46e-19
C12076 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 2.33e-19
C12077 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00594f
C12078 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# sky130_fd_sc_hd__inv_1_105/Y 6.69e-19
C12079 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 6.64e-20
C12080 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.72e-20
C12081 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 0.00944f
C12082 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__inv_1_18/Y 0.00357f
C12083 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__inv_1_9/Y 0.00127f
C12084 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__conb_1_5/HI 2.15e-20
C12085 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 2.75e-20
C12086 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# V_LOW 0.00706f
C12087 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_42/HI 0.107f
C12088 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__nand2_8_9/Y 3.21e-20
C12089 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0109f
C12090 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# V_LOW 0.0353f
C12091 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_27_47# 0.07f
C12092 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# sky130_fd_sc_hd__conb_1_26/HI -2.65e-20
C12093 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_16/LO 5.37e-21
C12094 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 9.11e-21
C12095 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00206f
C12096 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# V_LOW 0.00377f
C12097 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0413f
C12098 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0395f
C12099 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -7.6e-19
C12100 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# -5.54e-21
C12101 FULL_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 2.43f
C12102 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 6.83e-20
C12103 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# sky130_fd_sc_hd__inv_1_18/Y 1.69e-19
C12104 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.42e-19
C12105 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__conb_1_47/HI 2.27e-21
C12106 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_19/Q_N 2.08e-21
C12107 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# sky130_fd_sc_hd__conb_1_6/HI -1.25e-20
C12108 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0107f
C12109 FULL_COUNTER.COUNT_SUB_DFF12.Q V_GND 2.8f
C12110 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 1.33e-19
C12111 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00707f
C12112 FULL_COUNTER.COUNT_SUB_DFF10.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 1.27f
C12113 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00221f
C12114 sky130_fd_sc_hd__inv_1_109/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.127f
C12115 sky130_fd_sc_hd__inv_1_97/Y sky130_fd_sc_hd__inv_1_93/A 2.74e-19
C12116 RISING_COUNTER.COUNT_SUB_DFF11.Q V_GND 1.37f
C12117 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# V_LOW 1.38e-19
C12118 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__inv_1_57/Y 0.0157f
C12119 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 6.15e-19
C12120 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# V_GND 4.69e-19
C12121 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 0.0398f
C12122 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00649f
C12123 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# V_GND 0.00395f
C12124 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__inv_1_99/Y 0.0669f
C12125 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# V_LOW 0.0222f
C12126 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.46e-19
C12127 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0245f
C12128 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0193f
C12129 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_72/A 7.93e-20
C12130 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# V_LOW 0.0198f
C12131 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# V_GND 0.00646f
C12132 sky130_fd_sc_hd__dfbbn_1_43/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 9.68e-20
C12133 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_75/A 6.36e-19
C12134 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# sky130_fd_sc_hd__conb_1_21/HI 1.26e-19
C12135 sky130_fd_sc_hd__conb_1_27/HI RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00241f
C12136 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__conb_1_40/HI 0.0173f
C12137 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 5.49e-20
C12138 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.00589f
C12139 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 1.08e-19
C12140 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 1.13e-19
C12141 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0.0072f
C12142 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 9.04e-20
C12143 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_581_47# -2.6e-20
C12144 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# -7.5e-20
C12145 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# sky130_fd_sc_hd__inv_1_6/Y 7.97e-21
C12146 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_1_107/Y 0.00846f
C12147 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_17/HI 6.55e-19
C12148 sky130_fd_sc_hd__dfbbn_1_22/a_581_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.96e-19
C12149 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.32e-19
C12150 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# sky130_fd_sc_hd__inv_1_98/Y 3.94e-21
C12151 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_12/Y 5.97e-20
C12152 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# V_GND 0.00102f
C12153 sky130_fd_sc_hd__nand3_1_0/Y V_LOW 0.514f
C12154 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 5.44e-19
C12155 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.05e-20
C12156 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# V_GND 3.32e-19
C12157 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# V_LOW 0.00685f
C12158 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__conb_1_38/HI 0.0206f
C12159 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_105/Y 0.187f
C12160 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_1_13/Y 1.97e-21
C12161 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.37e-22
C12162 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# V_GND 2.18e-19
C12163 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00131f
C12164 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# V_LOW 0.00163f
C12165 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.4e-21
C12166 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_39/LO 8.84e-20
C12167 sky130_fd_sc_hd__inv_1_51/A V_LOW 0.26f
C12168 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 4.72e-19
C12169 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_1_98/Y 0.00884f
C12170 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# -1.46e-19
C12171 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# -0.00183f
C12172 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# -4.1e-19
C12173 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_891_329# -2.2e-20
C12174 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_1_101/Y 3.09e-20
C12175 Reset sky130_fd_sc_hd__inv_1_119/Y 0.885f
C12176 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 0.0142f
C12177 sky130_fd_sc_hd__inv_1_17/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 1.11e-19
C12178 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 2.45e-20
C12179 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 2.4e-20
C12180 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 9.07e-21
C12181 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 8.8e-22
C12182 sky130_fd_sc_hd__nand2_8_2/A V_LOW 0.0454f
C12183 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# sky130_fd_sc_hd__conb_1_30/HI -2.07e-19
C12184 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_93/A 0.0026f
C12185 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 6.01e-21
C12186 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__conb_1_26/HI 1.86e-19
C12187 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# -2.74e-21
C12188 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -2.18e-19
C12189 sky130_fd_sc_hd__dfbbn_1_21/Q_N V_LOW -0.00509f
C12190 sky130_fd_sc_hd__dfbbn_1_47/Q_N CLOCK_GEN.SR_Op.Q 0.016f
C12191 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# V_LOW -0.108f
C12192 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.21e-19
C12193 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# 0.0019f
C12194 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__conb_1_35/HI 5.79e-19
C12195 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 9.59e-22
C12196 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 4.37e-20
C12197 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# V_GND -0.0105f
C12198 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 2.15e-19
C12199 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# sky130_fd_sc_hd__conb_1_22/HI 0.0024f
C12200 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# V_GND -0.00797f
C12201 sky130_fd_sc_hd__dfbbn_1_4/Q_N FULL_COUNTER.COUNT_SUB_DFF10.Q 4.09e-20
C12202 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# -0.00734f
C12203 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_891_329# -0.00159f
C12204 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__conb_1_34/LO 2.1e-19
C12205 sky130_fd_sc_hd__nand2_1_5/a_113_47# V_GND 4.29e-20
C12206 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.02e-19
C12207 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 7.08e-21
C12208 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__inv_1_9/Y 0.00207f
C12209 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.7e-20
C12210 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_27/Y 5.16e-20
C12211 sky130_fd_sc_hd__inv_1_55/Y sky130_fd_sc_hd__conb_1_30/HI 9.19e-19
C12212 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.0132f
C12213 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_63/Y 3.58e-20
C12214 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# V_LOW 4.5e-19
C12215 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00592f
C12216 sky130_fd_sc_hd__dfbbn_1_42/a_1340_413# V_LOW 2.94e-20
C12217 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.0448f
C12218 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_40/HI 0.0331f
C12219 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0588f
C12220 sky130_fd_sc_hd__dfbbn_1_8/Q_N FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0197f
C12221 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0553f
C12222 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 4.06e-21
C12223 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 2.07e-20
C12224 sky130_fd_sc_hd__conb_1_2/LO FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00942f
C12225 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.12e-19
C12226 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00547f
C12227 sky130_fd_sc_hd__inv_1_63/Y V_GND 0.0974f
C12228 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# V_GND -0.00506f
C12229 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.82e-19
C12230 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_66/Y 6.17e-20
C12231 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF0.Q 1e-20
C12232 sky130_fd_sc_hd__dfbbn_1_38/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 2.26e-19
C12233 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 8.9e-19
C12234 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 3.79e-20
C12235 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__conb_1_39/HI -0.00833f
C12236 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.81e-19
C12237 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# CLOCK_GEN.SR_Op.Q 2.15e-19
C12238 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 1.22e-19
C12239 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_43/Y 0.00101f
C12240 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.15e-20
C12241 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__inv_1_18/Y 0.0141f
C12242 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_4/Y 0.0172f
C12243 sky130_fd_sc_hd__inv_1_95/A V_GND 0.484f
C12244 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00466f
C12245 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_20/Y 0.00144f
C12246 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_891_329# -2.2e-20
C12247 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# -0.00459f
C12248 sky130_fd_sc_hd__dfbbn_1_21/a_581_47# sky130_fd_sc_hd__inv_1_57/Y 3.73e-19
C12249 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__conb_1_18/HI 4.1e-19
C12250 sky130_fd_sc_hd__nand3_1_1/a_109_47# V_GND 1.15e-19
C12251 sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# sky130_fd_sc_hd__inv_16_1/Y 0.00485f
C12252 sky130_fd_sc_hd__dfbbn_1_42/a_1159_47# V_GND 8.06e-19
C12253 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_473_413# -0.012f
C12254 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -0.00701f
C12255 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# V_LOW -0.00423f
C12256 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0355f
C12257 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.83e-19
C12258 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_32/HI 0.0213f
C12259 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# sky130_fd_sc_hd__conb_1_35/HI 2.63e-19
C12260 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# V_LOW 0.00508f
C12261 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# V_GND 0.00689f
C12262 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__conb_1_21/HI 2.95e-19
C12263 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.15e-19
C12264 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# -1.24e-20
C12265 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# Reset 8.41e-19
C12266 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 4.87e-20
C12267 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.08e-20
C12268 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 2.02e-22
C12269 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 9.45e-21
C12270 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 5.19e-19
C12271 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 1.97e-19
C12272 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/Q_N -4.33e-20
C12273 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0129f
C12274 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.26e-37
C12275 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.52e-21
C12276 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q -4.98e-20
C12277 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_8/HI 0.0155f
C12278 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_23/Y 2.37e-20
C12279 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# sky130_fd_sc_hd__nand3_1_0/Y 2.02e-19
C12280 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__inv_1_4/Y 9.79e-21
C12281 sky130_fd_sc_hd__dfbbn_1_49/a_1340_413# sky130_fd_sc_hd__conb_1_38/HI 4.53e-19
C12282 sky130_fd_sc_hd__dfbbn_1_45/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 6e-20
C12283 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_53/Y 3.01e-19
C12284 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_22/HI 1.35e-19
C12285 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 3.68e-19
C12286 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# sky130_fd_sc_hd__conb_1_28/HI -4.57e-19
C12287 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__conb_1_9/LO 9.06e-20
C12288 sky130_fd_sc_hd__inv_1_62/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 1.49e-21
C12289 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.43e-21
C12290 sky130_fd_sc_hd__dfbbn_1_20/a_557_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.03e-19
C12291 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__inv_1_98/Y 0.0374f
C12292 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# -7.47e-20
C12293 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 7.58e-20
C12294 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# 1.42e-32
C12295 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# -0.00385f
C12296 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 4.65e-20
C12297 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 2.74e-21
C12298 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 5.95e-21
C12299 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__conb_1_17/HI 5.06e-20
C12300 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -0.00932f
C12301 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_473_413# -0.012f
C12302 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__conb_1_17/HI 2.38e-19
C12303 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# -3.34e-20
C12304 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# V_LOW -9.94e-19
C12305 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00187f
C12306 RISING_COUNTER.COUNT_SUB_DFF14.Q V_GND 0.829f
C12307 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 8.26e-20
C12308 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# V_GND -0.0135f
C12309 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.33e-19
C12310 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# V_GND -0.00111f
C12311 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# -0.00592f
C12312 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_55/Y 0.0675f
C12313 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__inv_1_66/Y 8.49e-19
C12314 sky130_fd_sc_hd__conb_1_32/LO sky130_fd_sc_hd__conb_1_32/HI 0.0176f
C12315 sky130_fd_sc_hd__dfbbn_1_37/Q_N V_LOW 9.89e-19
C12316 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# V_LOW 0.00245f
C12317 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 1.81e-20
C12318 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# V_LOW 0.0102f
C12319 sky130_fd_sc_hd__conb_1_15/LO V_GND -0.00375f
C12320 sky130_fd_sc_hd__nand3_1_0/a_193_47# V_GND -9.68e-19
C12321 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_891_329# -2.2e-20
C12322 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# -0.00398f
C12323 sky130_fd_sc_hd__nand3_1_1/a_109_47# sky130_fd_sc_hd__nand3_1_1/Y 7.74e-19
C12324 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 0.00267f
C12325 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# sky130_fd_sc_hd__conb_1_40/HI 2.25e-19
C12326 sky130_fd_sc_hd__conb_1_46/LO sky130_fd_sc_hd__conb_1_49/HI 0.00288f
C12327 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/Q_N -4.78e-20
C12328 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 4.43e-21
C12329 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0127f
C12330 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_473_413# 0.00132f
C12331 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_14/Y 0.347f
C12332 sky130_fd_sc_hd__dfbbn_1_0/a_1363_47# V_GND -2.81e-19
C12333 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0306f
C12334 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 3.78e-19
C12335 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 3.29e-19
C12336 sky130_fd_sc_hd__dfbbn_1_20/a_581_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.02e-19
C12337 FULL_COUNTER.COUNT_SUB_DFF18.Q sky130_fd_sc_hd__conb_1_17/HI 0.405f
C12338 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__conb_1_39/HI -9.71e-19
C12339 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_26/HI 9.92e-19
C12340 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0103f
C12341 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.98e-21
C12342 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_100/Y 0.00575f
C12343 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.67e-19
C12344 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# -0.00552f
C12345 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 0.558f
C12346 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 2.83e-19
C12347 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# V_GND 0.00303f
C12348 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# V_GND 0.00205f
C12349 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# -2.57e-20
C12350 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# V_LOW 0.0138f
C12351 sky130_fd_sc_hd__dfbbn_1_22/a_1340_413# sky130_fd_sc_hd__conb_1_32/HI 5.29e-19
C12352 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0206f
C12353 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# sky130_fd_sc_hd__inv_1_112/Y 0.0072f
C12354 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0136f
C12355 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_581_47# -2.6e-20
C12356 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 1.75e-20
C12357 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__inv_1_78/A 6.97e-20
C12358 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_45/HI 0.0222f
C12359 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 9.4e-21
C12360 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.00459f
C12361 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0109f
C12362 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.13e-19
C12363 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_70/Y 0.00379f
C12364 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# sky130_fd_sc_hd__inv_1_5/Y 4.19e-19
C12365 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__nand2_1_0/Y 0.00375f
C12366 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.36e-20
C12367 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# -6.23e-21
C12368 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# -0.00149f
C12369 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_60/Y 0.00532f
C12370 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# Reset 0.00364f
C12371 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 8.11e-19
C12372 FALLING_COUNTER.COUNT_SUB_DFF11.Q FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0534f
C12373 sky130_fd_sc_hd__conb_1_23/HI V_LOW 0.00899f
C12374 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# V_GND 0.00176f
C12375 sky130_fd_sc_hd__inv_1_98/Y Reset 0.0416f
C12376 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00259f
C12377 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.204f
C12378 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_94/A 0.134f
C12379 sky130_fd_sc_hd__conb_1_25/HI V_LOW 0.0831f
C12380 RISING_COUNTER.COUNT_SUB_DFF12.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0411f
C12381 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 2.54e-20
C12382 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 5.08e-20
C12383 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__inv_1_90/Y 5.04e-20
C12384 sky130_fd_sc_hd__nand2_1_3/a_113_47# V_GND 3.2e-20
C12385 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__conb_1_11/HI 7.88e-22
C12386 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_2/a_27_47# 7.23e-20
C12387 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_30/LO 5.12e-20
C12388 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 1e-19
C12389 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/Q_N -4.33e-20
C12390 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.62e-20
C12391 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_473_413# -0.0144f
C12392 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_647_21# -0.0105f
C12393 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 4.14e-20
C12394 sky130_fd_sc_hd__inv_1_111/Y V_GND 0.0361f
C12395 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# CLOCK_GEN.SR_Op.Q 5.81e-21
C12396 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_32/a_1340_413# -2.57e-20
C12397 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 2.11e-19
C12398 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__conb_1_17/HI 4.32e-20
C12399 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__conb_1_9/HI 2.08e-21
C12400 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/Q_N -4.24e-20
C12401 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.92e-21
C12402 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 1.81e-20
C12403 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/Q_N -6.48e-19
C12404 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 3.29e-19
C12405 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# V_LOW 0.00185f
C12406 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# -5.54e-21
C12407 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# -0.00138f
C12408 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_112/Y 0.00941f
C12409 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.66e-20
C12410 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_1159_47# 1.2e-19
C12411 sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# V_LOW 1.79e-20
C12412 sky130_fd_sc_hd__fill_4_72/VPB V_LOW 0.797f
C12413 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# 1.42e-32
C12414 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# -0.00282f
C12415 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# sky130_fd_sc_hd__inv_1_57/Y 0.00134f
C12416 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 7.17e-21
C12417 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_97/Y 0.0281f
C12418 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_80/A 0.018f
C12419 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 3.25e-20
C12420 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# sky130_fd_sc_hd__inv_16_1/Y 1.38e-20
C12421 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 2.31e-20
C12422 sky130_fd_sc_hd__nand2_1_3/Y sky130_fd_sc_hd__inv_1_76/A 4.94e-19
C12423 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 1.2e-19
C12424 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.55e-19
C12425 sky130_fd_sc_hd__dfbbn_1_31/Q_N FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00232f
C12426 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_24/LO 3.47e-21
C12427 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.64e-19
C12428 sky130_fd_sc_hd__conb_1_19/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0106f
C12429 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0.0119f
C12430 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 0.00267f
C12431 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 9.59e-19
C12432 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 1.09e-19
C12433 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__conb_1_39/HI -2.17e-19
C12434 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__inv_1_102/Y 8.92e-19
C12435 sky130_fd_sc_hd__conb_1_0/HI sky130_fd_sc_hd__inv_16_2/Y 0.00168f
C12436 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00145f
C12437 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0.0383f
C12438 sky130_fd_sc_hd__conb_1_35/HI V_GND 0.0721f
C12439 sky130_fd_sc_hd__fill_4_69/VPB V_GND 0.4f
C12440 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# V_LOW 0.00729f
C12441 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_26/HI 6.56e-20
C12442 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.98e-20
C12443 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__conb_1_2/HI 0.00366f
C12444 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__conb_1_4/HI 0.032f
C12445 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_42/Y 0.0443f
C12446 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_1_98/Y 1.01e-21
C12447 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 2.41e-19
C12448 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.00893f
C12449 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# V_GND 0.00785f
C12450 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.82e-19
C12451 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# V_GND -0.00592f
C12452 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 1.11e-19
C12453 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# V_GND 1.74e-19
C12454 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0144f
C12455 sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# V_LOW 1.79e-20
C12456 RISING_COUNTER.COUNT_SUB_DFF0.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 5.56e-20
C12457 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_557_413# 1.25e-19
C12458 sky130_fd_sc_hd__dfbbn_1_41/a_1159_47# sky130_fd_sc_hd__inv_1_112/Y 5.98e-19
C12459 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00175f
C12460 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__inv_1_107/Y 0.0161f
C12461 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_1_99/Y 7.12e-20
C12462 sky130_fd_sc_hd__dfbbn_1_49/a_1112_329# sky130_fd_sc_hd__nand3_1_2/Y 1.1e-20
C12463 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.62e-21
C12464 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 5.71e-20
C12465 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# V_GND -0.183f
C12466 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.21e-20
C12467 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0.00103f
C12468 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__conb_1_0/HI 0.0143f
C12469 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# sky130_fd_sc_hd__inv_1_5/Y 4.31e-19
C12470 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# V_GND -0.00487f
C12471 sky130_fd_sc_hd__conb_1_20/LO CLOCK_GEN.SR_Op.Q 4.91e-19
C12472 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__conb_1_36/HI 0.0135f
C12473 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__inv_1_103/Y 0.0056f
C12474 sky130_fd_sc_hd__inv_1_105/Y V_LOW 0.256f
C12475 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00622f
C12476 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_791_47# 4.46e-20
C12477 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__inv_1_61/Y 1.07e-20
C12478 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_1_61/Y 1.63e-20
C12479 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__conb_1_11/HI 3.28e-19
C12480 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__conb_1_6/LO 1.06e-19
C12481 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# V_GND -3.53e-19
C12482 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# sky130_fd_sc_hd__conb_1_34/HI 2.1e-19
C12483 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.55e-19
C12484 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0312f
C12485 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_42/HI 0.0216f
C12486 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.7e-21
C12487 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__conb_1_45/HI 0.00537f
C12488 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__conb_1_38/HI 2.59e-19
C12489 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.15e-19
C12490 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# CLOCK_GEN.SR_Op.Q 4.06e-21
C12491 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__conb_1_24/HI 2.71e-19
C12492 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.45e-19
C12493 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.0404f
C12494 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.01f
C12495 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.0209f
C12496 sky130_fd_sc_hd__dfbbn_1_35/a_581_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 4.04e-20
C12497 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__conb_1_2/HI 0.00129f
C12498 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 5.11e-20
C12499 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# -0.00631f
C12500 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# -0.0147f
C12501 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 2.09e-21
C12502 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__inv_1_102/Y 0.0283f
C12503 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.3e-20
C12504 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0.0124f
C12505 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_108/Y 1.82e-19
C12506 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_1_4/Y 0.00373f
C12507 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 1.41e-20
C12508 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00165f
C12509 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_5/HI 0.117f
C12510 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_23/Y 0.0441f
C12511 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 9.08e-20
C12512 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__inv_1_75/A 0.00962f
C12513 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_65/Y 2.72e-19
C12514 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# -9.32e-20
C12515 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00455f
C12516 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.14e-20
C12517 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.64e-20
C12518 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__inv_1_15/Y 6.3e-19
C12519 FULL_COUNTER.COUNT_SUB_DFF3.Q V_LOW 5.92f
C12520 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 4.23e-21
C12521 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__conb_1_18/HI 2.98e-20
C12522 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 0.0123f
C12523 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# sky130_fd_sc_hd__conb_1_5/HI 1.21e-19
C12524 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_13/HI 0.00947f
C12525 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# 3.93e-19
C12526 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# V_LOW -9.15e-19
C12527 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 0.00222f
C12528 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 4.81e-20
C12529 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 3.89e-19
C12530 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.98e-19
C12531 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__conb_1_42/HI 0.0268f
C12532 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# sky130_fd_sc_hd__conb_1_2/HI 0.0063f
C12533 sky130_fd_sc_hd__inv_1_26/Y V_GND 0.117f
C12534 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__conb_1_4/HI 5.96e-19
C12535 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__nand2_8_0/a_27_47# 7.56e-19
C12536 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__inv_16_2/Y 3.63e-19
C12537 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_1_100/Y 5.61e-19
C12538 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__inv_1_98/Y 5.66e-21
C12539 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 7.19e-19
C12540 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_791_47# 9.78e-19
C12541 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 8.12e-19
C12542 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# V_GND 0.0202f
C12543 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_16_2/Y 4.43e-21
C12544 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_18/LO 2.86e-20
C12545 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# 6.85e-20
C12546 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF12.Q 0.249f
C12547 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__inv_1_58/Y 1.42e-19
C12548 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.022f
C12549 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# sky130_fd_sc_hd__inv_1_107/Y 8.57e-21
C12550 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_647_21# 0.00258f
C12551 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.121f
C12552 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.005f
C12553 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_10/HI 0.0152f
C12554 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0338f
C12555 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.59e-20
C12556 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_557_413# 9.73e-19
C12557 sky130_fd_sc_hd__dfbbn_1_10/a_1340_413# V_GND 1.13e-19
C12558 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_647_21# -6.43e-20
C12559 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# -5.78e-20
C12560 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__conb_1_10/HI 0.00159f
C12561 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# sky130_fd_sc_hd__conb_1_1/HI 0.00107f
C12562 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__conb_1_36/HI 0.01f
C12563 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# sky130_fd_sc_hd__conb_1_0/HI 6.43e-20
C12564 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# V_GND -0.00536f
C12565 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__inv_16_1/Y 6.54e-19
C12566 sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# sky130_fd_sc_hd__inv_1_103/Y 1.44e-21
C12567 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_94/Y 0.00216f
C12568 sky130_fd_sc_hd__dfbbn_1_39/a_581_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00242f
C12569 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 0.101f
C12570 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__conb_1_2/HI 0.0116f
C12571 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.03f
C12572 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# sky130_fd_sc_hd__conb_1_11/HI 0.00119f
C12573 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_51/HI 3.23e-20
C12574 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# V_GND 0.0251f
C12575 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_8_9/Y 4.03e-21
C12576 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.46e-20
C12577 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_19/Y 0.193f
C12578 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.0155f
C12579 sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# sky130_fd_sc_hd__conb_1_45/HI 2e-19
C12580 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__conb_1_38/HI 6.32e-19
C12581 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# V_GND -0.00113f
C12582 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_10/Y 0.0709f
C12583 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# sky130_fd_sc_hd__conb_1_24/HI 0.00198f
C12584 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# 0.00477f
C12585 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 6.63e-19
C12586 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 4.43e-21
C12587 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 0.0355f
C12588 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_35/LO 8.84e-20
C12589 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__conb_1_11/HI 6.27e-19
C12590 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__conb_1_45/LO 0.00434f
C12591 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00248f
C12592 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.79e-20
C12593 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_20/Y 1.31e-20
C12594 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# V_GND 0.00877f
C12595 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.95e-21
C12596 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_62/Y 0.00426f
C12597 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00105f
C12598 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# V_GND 8.51e-19
C12599 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__inv_1_21/Y 3.67e-19
C12600 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__nor2_1_0/Y 4.02e-20
C12601 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# sky130_fd_sc_hd__inv_1_4/Y 1.07e-21
C12602 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/Q_N -4.24e-20
C12603 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 0.0303f
C12604 sky130_fd_sc_hd__dfbbn_1_48/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.23e-19
C12605 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__inv_1_75/A 0.00501f
C12606 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF10.Q 1.16e-20
C12607 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.16f
C12608 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0123f
C12609 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.556f
C12610 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.02e-19
C12611 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__conb_1_43/LO 0.00126f
C12612 sky130_fd_sc_hd__fill_4_75/VPB V_GND 0.394f
C12613 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# -3.06e-20
C12614 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# -6.43e-20
C12615 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.39e-20
C12616 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# 0.00149f
C12617 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.89e-21
C12618 sky130_fd_sc_hd__dfbbn_1_19/a_1363_47# sky130_fd_sc_hd__conb_1_5/HI 3.38e-19
C12619 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 8.49e-22
C12620 sky130_fd_sc_hd__inv_1_103/Y sky130_fd_sc_hd__inv_16_1/Y 0.0237f
C12621 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_46/HI 3.36e-19
C12622 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.00996f
C12623 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 3.58e-19
C12624 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0974f
C12625 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__inv_1_100/Y 0.00134f
C12626 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# V_GND -0.00229f
C12627 sky130_fd_sc_hd__dfbbn_1_34/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00307f
C12628 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# -0.00216f
C12629 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_34/a_381_47# -0.00832f
C12630 sky130_fd_sc_hd__inv_1_6/Y Reset 1.03e-19
C12631 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__inv_1_22/Y 1.24e-19
C12632 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00555f
C12633 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 9.89e-19
C12634 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# V_LOW 3.56e-20
C12635 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00175f
C12636 sky130_fd_sc_hd__inv_1_88/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 0.168f
C12637 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# V_LOW 0.0158f
C12638 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__conb_1_27/HI 0.00196f
C12639 sky130_fd_sc_hd__conb_1_33/HI sky130_fd_sc_hd__nand3_1_0/Y 1.15e-19
C12640 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 9.23e-19
C12641 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.48e-21
C12642 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__inv_1_60/Y 0.00498f
C12643 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# V_LOW -0.109f
C12644 sky130_fd_sc_hd__dfbbn_1_6/a_581_47# sky130_fd_sc_hd__conb_1_10/HI 1.82e-19
C12645 Reset sky130_fd_sc_hd__nand2_1_0/Y 0.106f
C12646 sky130_fd_sc_hd__dfbbn_1_3/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.52e-19
C12647 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# V_LOW -0.00266f
C12648 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__conb_1_0/HI 1.38e-20
C12649 sky130_fd_sc_hd__dfbbn_1_32/Q_N V_GND -0.00787f
C12650 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__dfbbn_1_29/a_581_47# 3.72e-20
C12651 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 8.4e-19
C12652 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_47/HI -1.63e-20
C12653 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_381_47# 2.51e-19
C12654 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.08e-19
C12655 sky130_fd_sc_hd__inv_1_52/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 2.89e-20
C12656 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 1.31e-19
C12657 FULL_COUNTER.COUNT_SUB_DFF5.Q V_LOW 4.93f
C12658 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__conb_1_51/HI 5.86e-21
C12659 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__inv_1_61/Y 5.85e-22
C12660 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# V_LOW 4.8e-20
C12661 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 0.00149f
C12662 sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# V_GND 4.09e-19
C12663 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# V_LOW -0.00389f
C12664 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# -8.23e-19
C12665 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# -3.04e-19
C12666 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# V_GND -0.00424f
C12667 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# V_LOW 2.26e-20
C12668 sky130_fd_sc_hd__dfbbn_1_10/Q_N FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0247f
C12669 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_13/HI 1.62e-19
C12670 sky130_fd_sc_hd__nand2_8_2/A sky130_fd_sc_hd__inv_1_80/A 0.0199f
C12671 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_193_47# -0.154f
C12672 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 1.85e-19
C12673 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# V_GND -0.00521f
C12674 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0.00131f
C12675 sky130_fd_sc_hd__dfbbn_1_34/a_581_47# V_GND -8.97e-19
C12676 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# sky130_fd_sc_hd__conb_1_13/HI 1.49e-19
C12677 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_941_21# -1.62e-20
C12678 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# -2.41e-19
C12679 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0642f
C12680 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# V_LOW 0.00592f
C12681 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__conb_1_37/HI 0.00323f
C12682 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__conb_1_35/HI 0.00425f
C12683 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_1_107/Y 5.35e-19
C12684 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# V_GND 0.00347f
C12685 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 3.34e-19
C12686 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__conb_1_29/LO 0.00118f
C12687 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 3.05e-19
C12688 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 3.79e-19
C12689 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0.0095f
C12690 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 9.7e-20
C12691 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_941_21# -0.0597f
C12692 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00149f
C12693 sky130_fd_sc_hd__dfbbn_1_29/a_581_47# V_GND 4.43e-19
C12694 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# V_GND 7.54e-19
C12695 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# V_LOW 0.00658f
C12696 sky130_fd_sc_hd__inv_1_47/Y V_GND 0.121f
C12697 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.87e-20
C12698 sky130_fd_sc_hd__conb_1_0/HI sky130_fd_sc_hd__inv_1_9/Y 6.85e-19
C12699 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# V_LOW -0.0203f
C12700 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 0.0196f
C12701 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 3.07e-19
C12702 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# V_GND -0.00364f
C12703 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_85/A 0.0278f
C12704 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# V_LOW -0.115f
C12705 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.3e-19
C12706 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0264f
C12707 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.74e-19
C12708 sky130_fd_sc_hd__inv_1_71/Y V_LOW 0.251f
C12709 sky130_fd_sc_hd__conb_1_14/LO V_LOW 0.0556f
C12710 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 8.45e-21
C12711 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# V_GND 0.00456f
C12712 sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# V_LOW -0.00266f
C12713 sky130_fd_sc_hd__conb_1_18/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 0.234f
C12714 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# sky130_fd_sc_hd__conb_1_35/HI 1.11e-21
C12715 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0129f
C12716 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 0.00163f
C12717 sky130_fd_sc_hd__conb_1_40/HI sky130_fd_sc_hd__inv_16_1/Y 0.1f
C12718 sky130_fd_sc_hd__inv_1_110/Y FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.275f
C12719 sky130_fd_sc_hd__conb_1_16/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00518f
C12720 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 0.00668f
C12721 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.27e-20
C12722 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_647_21# -0.00791f
C12723 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 1.16e-21
C12724 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# Reset 0.00704f
C12725 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_62/Y 1.15e-20
C12726 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 4.58e-19
C12727 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_791_47# 7.44e-21
C12728 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 2.38e-20
C12729 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# V_GND -0.00404f
C12730 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_21/Y 0.00155f
C12731 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_20/Y 5.46e-20
C12732 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0.106f
C12733 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# V_GND 0.00335f
C12734 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00595f
C12735 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# -2.14e-19
C12736 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# V_GND 0.00183f
C12737 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__conb_1_27/LO 4.01e-19
C12738 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.324f
C12739 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# V_LOW -7.15e-19
C12740 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.67e-19
C12741 sky130_fd_sc_hd__dfbbn_1_36/a_581_47# V_GND -9.12e-19
C12742 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_25/LO 9.03e-20
C12743 RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_60/Y 5.16e-20
C12744 sky130_fd_sc_hd__inv_1_119/Y V_HIGH 0.435f
C12745 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0048f
C12746 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 8.75e-21
C12747 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.135f
C12748 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 7.78e-20
C12749 sky130_fd_sc_hd__dfbbn_1_20/a_581_47# V_LOW 9.05e-20
C12750 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__inv_1_13/Y 3.61e-21
C12751 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00635f
C12752 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_27/HI -2.07e-19
C12753 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_2/Y 2.24e-20
C12754 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.39e-21
C12755 sky130_fd_sc_hd__nand2_8_1/a_27_47# V_LOW -0.00847f
C12756 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__inv_1_21/Y 1.17e-19
C12757 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# V_LOW -9.94e-19
C12758 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# -0.00832f
C12759 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# -0.00242f
C12760 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# -6.22e-19
C12761 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 7.99e-19
C12762 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 7.99e-19
C12763 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__conb_1_44/LO 4.01e-19
C12764 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_44/HI 0.413f
C12765 sky130_fd_sc_hd__inv_1_15/Y V_LOW 0.121f
C12766 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# V_LOW -0.00266f
C12767 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# V_LOW 0.0162f
C12768 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__conb_1_47/HI -2.07e-19
C12769 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# V_GND 0.0159f
C12770 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__conb_1_46/HI 0.00422f
C12771 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_67/Y 0.259f
C12772 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 0.0287f
C12773 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0076f
C12774 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__inv_1_12/Y 0.00177f
C12775 sky130_fd_sc_hd__nand2_8_9/a_27_47# V_LOW -0.00528f
C12776 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_65/Y 0.0299f
C12777 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__conb_1_13/HI 4.06e-20
C12778 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_61/Y 0.132f
C12779 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 8.9e-21
C12780 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__conb_1_13/LO 3.38e-20
C12781 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 2.7e-22
C12782 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 0.0016f
C12783 sky130_fd_sc_hd__inv_1_68/Y sky130_fd_sc_hd__inv_1_67/Y 0.00157f
C12784 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__inv_1_12/Y 1.2e-19
C12785 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# V_GND -0.00502f
C12786 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_24/HI 4.75e-19
C12787 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 0.0172f
C12788 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 6.92e-21
C12789 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 5.77e-21
C12790 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 3.79e-20
C12791 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# V_GND 1.4e-19
C12792 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 0.0447f
C12793 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# V_LOW 0.0123f
C12794 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# sky130_fd_sc_hd__inv_1_9/Y 3.57e-19
C12795 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__conb_1_21/HI 4.43e-20
C12796 sky130_fd_sc_hd__fill_4_68/VPB V_LOW 0.797f
C12797 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# -1.76e-19
C12798 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 2.52e-20
C12799 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# -0.00486f
C12800 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_891_329# -0.00161f
C12801 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# sky130_fd_sc_hd__conb_1_37/HI 2.26e-21
C12802 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 8.6e-21
C12803 Reset RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0606f
C12804 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 1.13e-20
C12805 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# sky130_fd_sc_hd__conb_1_32/HI 0.0251f
C12806 sky130_fd_sc_hd__dfbbn_1_1/a_581_47# V_GND 1.97e-19
C12807 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00122f
C12808 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__inv_16_2/Y 8.69e-19
C12809 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# V_LOW 0.00249f
C12810 sky130_fd_sc_hd__dfbbn_1_9/a_557_413# V_GND 2.24e-19
C12811 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 2.44e-21
C12812 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_71/A 3.16e-20
C12813 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_16_1/Y 0.114f
C12814 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__inv_1_64/A 0.0244f
C12815 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_17/LO 0.0483f
C12816 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 3.6e-19
C12817 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__conb_1_13/HI 5.13e-19
C12818 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00246f
C12819 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__inv_1_22/Y 0.0501f
C12820 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_473_413# -3.86e-20
C12821 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -1.33e-19
C12822 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_15/LO 0.0141f
C12823 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0414f
C12824 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_891_329# 0.0017f
C12825 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.55e-20
C12826 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# V_LOW -7.17e-19
C12827 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__conb_1_44/HI -0.0119f
C12828 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 3.19e-19
C12829 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00217f
C12830 FULL_COUNTER.COUNT_SUB_DFF9.Q V_GND 1.1f
C12831 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# V_LOW -9.94e-19
C12832 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.99e-20
C12833 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# V_GND -0.0466f
C12834 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.45e-20
C12835 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 7.1e-19
C12836 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 6.33e-19
C12837 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.14e-19
C12838 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# V_GND 7.68e-19
C12839 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# Reset 0.0121f
C12840 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 1.85e-21
C12841 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 4.14e-21
C12842 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 8.79e-22
C12843 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 1.59e-19
C12844 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0507f
C12845 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00167f
C12846 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0.0019f
C12847 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# V_GND -0.00268f
C12848 sky130_fd_sc_hd__conb_1_51/LO FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0437f
C12849 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_24/HI 0.249f
C12850 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.872f
C12851 Reset sky130_fd_sc_hd__inv_1_65/Y 0.109f
C12852 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nand2_8_9/Y 0.00277f
C12853 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0184f
C12854 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_581_47# -2.6e-20
C12855 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# Reset 1.01e-19
C12856 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# sky130_fd_sc_hd__inv_1_62/Y 1.08e-20
C12857 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.7e-21
C12858 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0176f
C12859 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# 0.00423f
C12860 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.72e-19
C12861 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# V_GND 1.57e-19
C12862 sky130_fd_sc_hd__inv_1_53/Y V_GND 0.0317f
C12863 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_12/HI 0.0259f
C12864 sky130_fd_sc_hd__conb_1_30/LO V_LOW 0.0993f
C12865 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# -9.32e-20
C12866 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# -3.86e-20
C12867 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# -5.58e-20
C12868 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# V_GND 1.72e-19
C12869 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_98/Y 5.16e-20
C12870 sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__inv_16_0/Y 0.179f
C12871 sky130_fd_sc_hd__inv_1_55/Y RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0665f
C12872 sky130_fd_sc_hd__nand2_8_4/a_27_47# V_GND 0.054f
C12873 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# -4.84e-19
C12874 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# -5.54e-21
C12875 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 9.59e-19
C12876 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 0.00267f
C12877 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 0.0119f
C12878 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 1.09e-19
C12879 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.56e-21
C12880 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/Q_N -7.69e-20
C12881 FALLING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_108/Y 0.0735f
C12882 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 0.0879f
C12883 sky130_fd_sc_hd__dfbbn_1_21/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF2.Q 8.82e-19
C12884 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 1.42e-32
C12885 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -2.18e-19
C12886 FULL_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_1_12/Y 0.0339f
C12887 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 4.61e-20
C12888 sky130_fd_sc_hd__conb_1_41/LO V_LOW 0.0601f
C12889 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 2.53e-20
C12890 sky130_fd_sc_hd__conb_1_16/LO sky130_fd_sc_hd__inv_1_21/Y 8.37e-19
C12891 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# -0.00242f
C12892 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_381_47# -0.00201f
C12893 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 8.15e-20
C12894 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__conb_1_38/LO 5.4e-21
C12895 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 5.38e-19
C12896 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 8.75e-19
C12897 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 5.38e-19
C12898 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 8.75e-19
C12899 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 0.0107f
C12900 sky130_fd_sc_hd__conb_1_1/HI V_GND -0.131f
C12901 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 2.54e-20
C12902 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 7.07e-21
C12903 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 9.66e-19
C12904 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__conb_1_44/HI 9.6e-19
C12905 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 0.0124f
C12906 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__inv_1_102/Y 1.82e-19
C12907 FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0115f
C12908 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# sky130_fd_sc_hd__conb_1_47/HI 3.45e-19
C12909 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__dfbbn_1_38/a_647_21# 8.05e-20
C12910 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__conb_1_11/LO 0.00206f
C12911 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# V_LOW -1.46e-19
C12912 sky130_fd_sc_hd__conb_1_2/HI V_LOW 0.312f
C12913 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_36/HI 0.0175f
C12914 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__conb_1_46/HI 0.00188f
C12915 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# V_GND 0.00298f
C12916 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# 5.98e-19
C12917 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__inv_1_15/Y 9.49e-20
C12918 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__conb_1_22/HI 1.32e-19
C12919 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_40/HI 1.11e-20
C12920 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_23/Y 0.281f
C12921 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_9/a_381_47# 3.35e-20
C12922 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 8.46e-21
C12923 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__inv_1_49/Y -1.12e-19
C12924 sky130_fd_sc_hd__inv_1_85/A sky130_fd_sc_hd__inv_1_83/Y 0.016f
C12925 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 1.44e-20
C12926 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/Q_N -9.56e-20
C12927 sky130_fd_sc_hd__dfbbn_1_14/a_1363_47# sky130_fd_sc_hd__inv_1_12/Y 3.37e-19
C12928 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.03e-20
C12929 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 1.2e-20
C12930 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 9.18e-20
C12931 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# V_LOW -0.00216f
C12932 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 2.44e-19
C12933 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__conb_1_39/HI 2.55e-20
C12934 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 7.13e-21
C12935 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__inv_1_58/Y 0.00317f
C12936 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_581_47# 2.17e-19
C12937 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 5.21e-20
C12938 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# sky130_fd_sc_hd__conb_1_41/HI 0.0114f
C12939 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# V_GND -0.184f
C12940 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_2_0/Y 2.15e-19
C12941 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# -0.00282f
C12942 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_1_13/Y 0.0102f
C12943 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 3.21e-21
C12944 sky130_fd_sc_hd__dfbbn_1_23/a_581_47# sky130_fd_sc_hd__conb_1_32/HI 2.47e-19
C12945 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0827f
C12946 sky130_fd_sc_hd__dfbbn_1_11/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF18.Q 1.61e-19
C12947 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 1.55e-20
C12948 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_15/Y 2.18e-19
C12949 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_50/Y 0.00331f
C12950 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 5.71e-19
C12951 FULL_COUNTER.COUNT_SUB_DFF11.Q V_GND 1.13f
C12952 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0.00408f
C12953 sky130_fd_sc_hd__conb_1_19/LO sky130_fd_sc_hd__inv_16_2/Y 0.0166f
C12954 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00643f
C12955 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__inv_1_15/Y 0.0166f
C12956 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_40/a_1340_413# -2.57e-20
C12957 RISING_COUNTER.COUNT_SUB_DFF2.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.351f
C12958 sky130_fd_sc_hd__nor2_1_0/Y Reset 0.176f
C12959 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_19/Y 9.87e-21
C12960 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 1.09e-19
C12961 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 1.6e-19
C12962 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__conb_1_36/LO 3.32e-20
C12963 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.78e-19
C12964 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.77e-19
C12965 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.3e-19
C12966 sky130_fd_sc_hd__dfbbn_1_13/a_891_329# V_GND 5.04e-19
C12967 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# -0.0222f
C12968 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# -0.00452f
C12969 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# V_LOW 0.0156f
C12970 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# V_GND 3.04e-19
C12971 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 8.81e-21
C12972 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 4.97e-20
C12973 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 5.11e-20
C12974 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 4.92e-20
C12975 sky130_fd_sc_hd__dfbbn_1_40/Q_N V_GND -0.00763f
C12976 sky130_fd_sc_hd__nand2_8_4/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 1.46e-19
C12977 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# Reset 0.00134f
C12978 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 7.55e-19
C12979 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0388f
C12980 sky130_fd_sc_hd__nor2_1_0/a_109_297# CLOCK_GEN.SR_Op.Q 1.29e-19
C12981 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.29e-21
C12982 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_891_329# 8.83e-20
C12983 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 2.51e-20
C12984 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# V_GND -0.00397f
C12985 sky130_fd_sc_hd__inv_1_103/Y V_LOW 0.163f
C12986 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 6.43e-20
C12987 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 4.25e-21
C12988 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 3.1e-20
C12989 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# -0.00336f
C12990 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0603f
C12991 sky130_fd_sc_hd__dfbbn_1_29/Q_N Reset 0.00105f
C12992 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0449f
C12993 sky130_fd_sc_hd__dfbbn_1_10/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 3.67e-20
C12994 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.00108f
C12995 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 4.99e-19
C12996 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 9.54e-19
C12997 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00418f
C12998 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0174f
C12999 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/Q_N -4.24e-20
C13000 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_6/a_1340_413# -2.57e-20
C13001 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 0.0174f
C13002 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# V_GND 0.00185f
C13003 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# sky130_fd_sc_hd__conb_1_51/HI 0.00173f
C13004 sky130_fd_sc_hd__inv_1_90/Y V_GND 0.0669f
C13005 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# -9.32e-20
C13006 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_1112_329# 2.07e-21
C13007 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__conb_1_37/HI 0.0116f
C13008 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 2.81e-20
C13009 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 4.35e-19
C13010 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# V_LOW 0.0205f
C13011 sky130_fd_sc_hd__nand2_1_2/A V_GND 0.122f
C13012 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_1340_413# 0.00148f
C13013 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.57e-20
C13014 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_381_47# 0.00453f
C13015 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 6.66e-21
C13016 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 2.19e-19
C13017 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__dfbbn_1_27/a_381_47# 2.19e-19
C13018 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# -3.34e-20
C13019 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_25/LO 0.0125f
C13020 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_16_2/Y 8.87e-19
C13021 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 0.00119f
C13022 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 7.15e-19
C13023 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 6.43e-19
C13024 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00378f
C13025 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/Q_N -9.56e-20
C13026 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# V_LOW -9.15e-19
C13027 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00715f
C13028 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_381_47# -0.00171f
C13029 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 5.96e-19
C13030 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# V_LOW 0.0264f
C13031 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# CLOCK_GEN.SR_Op.Q 6.44e-21
C13032 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__inv_1_13/Y 0.0135f
C13033 sky130_fd_sc_hd__dfbbn_1_4/Q_N V_GND 0.00173f
C13034 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__inv_1_8/Y 1.07e-20
C13035 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# V_LOW 1.38e-19
C13036 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# V_GND 0.00228f
C13037 sky130_fd_sc_hd__inv_1_16/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 1.2e-20
C13038 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__nand2_1_3/Y 0.0367f
C13039 sky130_fd_sc_hd__inv_1_27/Y V_SENSE 0.142f
C13040 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# 0.00158f
C13041 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.44e-19
C13042 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# V_LOW 3.93e-20
C13043 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 5.1e-19
C13044 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.21e-19
C13045 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/Q_N 1.54e-20
C13046 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__inv_1_9/Y 0.0314f
C13047 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# sky130_fd_sc_hd__conb_1_41/HI 0.0174f
C13048 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 4.74e-22
C13049 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 7.46e-21
C13050 sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# V_GND 1.06e-19
C13051 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__inv_1_90/Y 0.00132f
C13052 sky130_fd_sc_hd__inv_1_17/Y V_LOW 0.137f
C13053 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 0.002f
C13054 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0.00635f
C13055 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 9.18e-19
C13056 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/Q_N -6.48e-19
C13057 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_16_1/Y 0.284f
C13058 sky130_fd_sc_hd__dfbbn_1_44/Q_N sky130_fd_sc_hd__conb_1_26/LO 1.62e-20
C13059 FALLING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_40/HI 0.00712f
C13060 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__conb_1_13/HI 2.46e-20
C13061 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 7.56e-19
C13062 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_12/LO 0.0242f
C13063 sky130_fd_sc_hd__dfbbn_1_43/a_557_413# V_GND 2.37e-19
C13064 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__inv_1_15/Y 2.18e-19
C13065 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 7.41e-19
C13066 sky130_fd_sc_hd__dfbbn_1_3/a_1112_329# V_GND 0.00101f
C13067 sky130_fd_sc_hd__dfbbn_1_14/a_581_47# sky130_fd_sc_hd__inv_1_15/Y 6.57e-19
C13068 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 1.31e-19
C13069 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_55/Y 0.00493f
C13070 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 3.49e-19
C13071 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_1_16/Y 0.00362f
C13072 sky130_fd_sc_hd__dfbbn_1_34/a_557_413# sky130_fd_sc_hd__inv_1_103/Y 5.67e-19
C13073 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_23/Y 2.43e-20
C13074 sky130_fd_sc_hd__conb_1_4/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00895f
C13075 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__inv_1_23/Y 6.97e-21
C13076 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# -6.8e-19
C13077 sky130_fd_sc_hd__conb_1_40/HI V_LOW 0.141f
C13078 sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# V_LOW 1.79e-20
C13079 sky130_fd_sc_hd__conb_1_32/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 0.0413f
C13080 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 1.88e-19
C13081 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 1.6e-20
C13082 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 4.68e-20
C13083 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_473_413# -0.0222f
C13084 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -0.0133f
C13085 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 0.00329f
C13086 sky130_fd_sc_hd__dfbbn_1_1/Q_N Reset 0.00139f
C13087 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.00378f
C13088 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__conb_1_35/HI 0.021f
C13089 sky130_fd_sc_hd__dfbbn_1_14/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 2.98e-20
C13090 sky130_fd_sc_hd__conb_1_49/LO V_GND -0.00515f
C13091 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# Reset 5.77e-19
C13092 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.28e-21
C13093 sky130_fd_sc_hd__dfbbn_1_7/Q_N V_GND -0.00775f
C13094 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 2.87e-20
C13095 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__conb_1_45/HI 0.0246f
C13096 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 9.39e-20
C13097 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 0.00107f
C13098 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 2.23e-19
C13099 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 5.64e-20
C13100 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0123f
C13101 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 1.16e-19
C13102 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0134f
C13103 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.02e-20
C13104 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_75/Y 1.08e-19
C13105 sky130_fd_sc_hd__dfbbn_1_24/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00814f
C13106 sky130_fd_sc_hd__conb_1_49/LO sky130_fd_sc_hd__inv_1_106/Y 3.82e-19
C13107 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.084f
C13108 sky130_fd_sc_hd__dfbbn_1_49/a_1363_47# V_GND -3.69e-19
C13109 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/Q_N -4.33e-20
C13110 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.23e-19
C13111 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1_17/HI 1.47e-21
C13112 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 1.86e-20
C13113 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0.00134f
C13114 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 1.28e-20
C13115 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# V_LOW 1.79e-20
C13116 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00133f
C13117 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_1363_47# 5.86e-20
C13118 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/Q_N -4.24e-20
C13119 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 2.84e-20
C13120 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 8.66e-20
C13121 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00169f
C13122 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 9.87e-20
C13123 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 0.00171f
C13124 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00295f
C13125 sky130_fd_sc_hd__dfbbn_1_8/a_557_413# sky130_fd_sc_hd__inv_16_2/Y 1.16e-19
C13126 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 1.83e-20
C13127 sky130_fd_sc_hd__dfbbn_1_25/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 8.62e-20
C13128 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/Q_N -9.56e-20
C13129 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__conb_1_46/HI 0.00201f
C13130 sky130_fd_sc_hd__dfbbn_1_1/a_557_413# sky130_fd_sc_hd__conb_1_2/HI 2.63e-19
C13131 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_76/A 0.02f
C13132 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0354f
C13133 sky130_fd_sc_hd__inv_1_56/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 1.56e-21
C13134 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# -1.44e-20
C13135 sky130_fd_sc_hd__dfbbn_1_36/a_557_413# sky130_fd_sc_hd__inv_1_103/Y 5.21e-19
C13136 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__inv_1_15/Y 2.05e-19
C13137 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__inv_16_2/Y 4.03e-20
C13138 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 3.59e-21
C13139 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__conb_1_19/LO 3.17e-20
C13140 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 0.0105f
C13141 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# V_LOW 0.011f
C13142 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__conb_1_47/HI 0.00102f
C13143 FALLING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__conb_1_46/HI 1.1e-19
C13144 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__inv_1_15/Y 1.14e-21
C13145 sky130_fd_sc_hd__dfbbn_1_17/a_1363_47# V_GND 1.72e-19
C13146 sky130_fd_sc_hd__inv_2_0/Y V_LOW 0.558f
C13147 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 2.5e-19
C13148 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 3.33e-19
C13149 sky130_fd_sc_hd__nand2_8_7/a_27_47# V_GND 0.0482f
C13150 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_53/Y 0.0263f
C13151 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_27/Q_N 3.26e-19
C13152 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_891_329# 0.00102f
C13153 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 8.85e-19
C13154 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 5.14e-20
C13155 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 2.27e-20
C13156 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 3.34e-19
C13157 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__conb_1_45/HI 0.0471f
C13158 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 0.0207f
C13159 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 3.56e-19
C13160 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 3.82e-19
C13161 sky130_fd_sc_hd__dfbbn_1_13/Q_N V_LOW -0.00497f
C13162 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# V_LOW 0.0122f
C13163 sky130_fd_sc_hd__inv_1_58/Y sky130_fd_sc_hd__inv_1_57/Y 0.0483f
C13164 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 1.48e-20
C13165 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 4.34e-20
C13166 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# V_LOW 0.0302f
C13167 sky130_fd_sc_hd__dfbbn_1_30/Q_N sky130_fd_sc_hd__conb_1_41/HI 0.0384f
C13168 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 9.36e-21
C13169 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 9.05e-20
C13170 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 0.00116f
C13171 sky130_fd_sc_hd__conb_1_37/HI sky130_fd_sc_hd__inv_1_91/Y 1.2e-20
C13172 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF19.Q 0.171f
C13173 sky130_fd_sc_hd__inv_1_85/A V_LOW 0.52f
C13174 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.582f
C13175 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.558f
C13176 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# V_LOW -0.318f
C13177 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.02f
C13178 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 5.19e-20
C13179 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__inv_16_1/Y 0.00105f
C13180 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0136f
C13181 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.00421f
C13182 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_381_47# -3.79e-20
C13183 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__dfbbn_1_46/a_1112_329# -4.66e-20
C13184 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__inv_1_54/Y 7.52e-21
C13185 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 0.00183f
C13186 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 1.76e-19
C13187 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 0.00183f
C13188 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 1.76e-19
C13189 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# V_LOW 0.0211f
C13190 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_5/Y 0.00114f
C13191 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# V_GND -0.0466f
C13192 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# V_GND -0.00112f
C13193 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# sky130_fd_sc_hd__conb_1_22/HI 2.54e-20
C13194 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__inv_1_23/Y 0.0108f
C13195 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# -0.00152f
C13196 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 0.0295f
C13197 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 9.81e-19
C13198 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# V_GND 2.6e-19
C13199 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# V_GND 0.00397f
C13200 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# -5.14e-19
C13201 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 3.11e-20
C13202 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 7.03e-21
C13203 FALLING_COUNTER.COUNT_SUB_DFF6.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.49f
C13204 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# V_GND -0.0441f
C13205 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__conb_1_35/HI 2.62e-20
C13206 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# sky130_fd_sc_hd__conb_1_45/HI 3.53e-19
C13207 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 2.16e-20
C13208 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_47/LO 8.09e-21
C13209 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_8_3/Y 0.00392f
C13210 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 1.04e-19
C13211 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 3.96e-19
C13212 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.00161f
C13213 sky130_fd_sc_hd__fill_4_74/VPB V_LOW 0.797f
C13214 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 7.69e-19
C13215 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__conb_1_49/HI 5.94e-19
C13216 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0042f
C13217 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__inv_1_106/Y 4.93e-19
C13218 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# V_GND -0.0431f
C13219 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_78/A 0.0357f
C13220 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# V_GND 0.00948f
C13221 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# 3.44e-20
C13222 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0371f
C13223 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 3.73e-20
C13224 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00603f
C13225 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 3.61e-19
C13226 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 2.81e-19
C13227 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__inv_1_11/Y 1.51e-19
C13228 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__nand3_1_0/Y 7.79e-19
C13229 sky130_fd_sc_hd__dfbbn_1_17/a_581_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.99e-19
C13230 sky130_fd_sc_hd__inv_1_50/A V_GND 0.336f
C13231 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# V_LOW 0.0163f
C13232 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0593f
C13233 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# 4.05e-21
C13234 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_1_23/Y 0.00237f
C13235 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 1.92e-19
C13236 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 5.78e-19
C13237 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 3.85e-19
C13238 sky130_fd_sc_hd__conb_1_30/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00606f
C13239 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00514f
C13240 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__inv_1_20/Y 0.0349f
C13241 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_42/LO 0.0111f
C13242 sky130_fd_sc_hd__inv_1_70/Y V_LOW 0.391f
C13243 sky130_fd_sc_hd__conb_1_26/LO RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0545f
C13244 sky130_fd_sc_hd__dfbbn_1_29/a_1112_329# sky130_fd_sc_hd__conb_1_33/HI 0.00138f
C13245 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# sky130_fd_sc_hd__conb_1_46/HI -2.07e-19
C13246 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_76/A 1.73e-19
C13247 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_381_47# -3.79e-20
C13248 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# -4.66e-20
C13249 sky130_fd_sc_hd__inv_1_110/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.72e-19
C13250 sky130_fd_sc_hd__inv_1_100/Y sky130_fd_sc_hd__conb_1_35/HI 2.56e-21
C13251 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_12/HI 2.27e-20
C13252 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.99e-19
C13253 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__inv_1_21/Y 8.53e-19
C13254 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 9.1e-21
C13255 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.0426f
C13256 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__inv_1_20/Y 1.07e-20
C13257 sky130_fd_sc_hd__dfbbn_1_16/Q_N sky130_fd_sc_hd__inv_1_8/Y 5.85e-22
C13258 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.9e-21
C13259 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__conb_1_50/HI 0.00174f
C13260 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# -0.00631f
C13261 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# -0.0119f
C13262 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.444f
C13263 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# V_GND -0.0203f
C13264 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__inv_1_11/Y 0.0339f
C13265 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 1.85e-19
C13266 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 6.05e-19
C13267 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.81e-21
C13268 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 3.7e-22
C13269 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 6.85e-20
C13270 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 0.00907f
C13271 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# sky130_fd_sc_hd__conb_1_45/HI 5.98e-19
C13272 sky130_fd_sc_hd__dfbbn_1_26/a_1112_329# V_LOW -0.00266f
C13273 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_1340_413# 1.57e-19
C13274 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__inv_1_17/Y 8.36e-19
C13275 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.33e-20
C13276 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# 8.99e-20
C13277 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 1.07e-20
C13278 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# V_LOW 0.018f
C13279 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# V_LOW 4.8e-20
C13280 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 7.31e-19
C13281 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_1_9/Y 7.32e-20
C13282 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_891_329# -0.00159f
C13283 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# -0.0079f
C13284 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/Q_N 0.00106f
C13285 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_1_100/Y 5.32e-20
C13286 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00204f
C13287 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__conb_1_46/HI 1.9e-20
C13288 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 7.78e-20
C13289 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# 2.3e-19
C13290 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 3.33e-19
C13291 sky130_fd_sc_hd__inv_1_61/Y sky130_fd_sc_hd__conb_1_28/HI 7e-19
C13292 sky130_fd_sc_hd__conb_1_12/LO sky130_fd_sc_hd__conb_1_17/HI 7.36e-19
C13293 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 6.88e-20
C13294 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 3.75e-19
C13295 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 0.00944f
C13296 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0.00944f
C13297 sky130_fd_sc_hd__inv_1_93/Y sky130_fd_sc_hd__inv_1_93/A 0.00734f
C13298 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_17/Y 0.041f
C13299 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# V_GND 2.47e-19
C13300 sky130_fd_sc_hd__dfbbn_1_26/a_581_47# V_GND -9.06e-19
C13301 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# sky130_fd_sc_hd__conb_1_22/HI 4.98e-19
C13302 sky130_fd_sc_hd__dfbbn_1_44/a_891_329# V_LOW 2.26e-20
C13303 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_105/Y 0.113f
C13304 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_581_47# -2.6e-20
C13305 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__nand2_8_9/Y 7.24e-19
C13306 sky130_fd_sc_hd__dfbbn_1_4/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 2.02e-19
C13307 sky130_fd_sc_hd__dfbbn_1_31/a_581_47# V_GND 2.05e-19
C13308 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_40/A 0.0366f
C13309 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 6.47e-19
C13310 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 2.99e-19
C13311 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 6.9e-19
C13312 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# V_GND 2.56e-19
C13313 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# V_LOW 0.0247f
C13314 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 0.00113f
C13315 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# V_GND 0.00309f
C13316 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_891_329# -2.46e-19
C13317 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_557_413# -3.67e-20
C13318 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# -0.00467f
C13319 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# CLOCK_GEN.SR_Op.Q 4.15e-19
C13320 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__conb_1_38/HI 0.0011f
C13321 sky130_fd_sc_hd__nand2_8_3/a_27_47# sky130_fd_sc_hd__nand2_1_5/Y 0.0104f
C13322 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0.00451f
C13323 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 8.46e-20
C13324 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__conb_1_11/HI 0.00102f
C13325 sky130_fd_sc_hd__nand3_1_2/B sky130_fd_sc_hd__inv_1_76/A 0.0205f
C13326 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 9.95e-20
C13327 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.72e-20
C13328 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0355f
C13329 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 5.58e-20
C13330 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_557_413# -3.67e-20
C13331 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_50/a_891_329# -2.46e-19
C13332 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# -0.0145f
C13333 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# 2.07e-21
C13334 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.9e-21
C13335 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# sky130_fd_sc_hd__conb_1_49/HI -2.86e-20
C13336 sky130_fd_sc_hd__dfbbn_1_23/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00904f
C13337 sky130_fd_sc_hd__conb_1_33/LO V_GND -0.00221f
C13338 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# sky130_fd_sc_hd__inv_1_106/Y 3.83e-19
C13339 sky130_fd_sc_hd__dfbbn_1_18/a_1672_329# V_GND 2.6e-19
C13340 sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# sky130_fd_sc_hd__inv_1_59/Y 6.65e-20
C13341 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# V_GND 0.00189f
C13342 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 4.01e-19
C13343 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 1.08e-20
C13344 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_42/HI 4.11e-19
C13345 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# Reset 0.00379f
C13346 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 8.63e-19
C13347 sky130_fd_sc_hd__dfbbn_1_19/a_557_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00269f
C13348 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 8.33e-19
C13349 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__inv_1_11/Y 2.89e-19
C13350 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.556f
C13351 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# -0.00864f
C13352 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# -0.0129f
C13353 sky130_fd_sc_hd__dfbbn_1_51/a_557_413# V_GND 2.42e-19
C13354 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.00361f
C13355 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0195f
C13356 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# 1.84e-21
C13357 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 5.71e-21
C13358 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# -2.18e-19
C13359 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# -5.54e-21
C13360 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.116f
C13361 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__inv_1_10/Y 0.00541f
C13362 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0457f
C13363 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.0078f
C13364 sky130_fd_sc_hd__dfbbn_1_5/Q_N FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0266f
C13365 sky130_fd_sc_hd__conb_1_22/LO RISING_COUNTER.COUNT_SUB_DFF11.Q 9.86e-21
C13366 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.0235f
C13367 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# -3.48e-20
C13368 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_891_329# -2.2e-20
C13369 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.43e-21
C13370 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 9.9e-20
C13371 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.56e-19
C13372 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__conb_1_2/HI 0.00856f
C13373 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 3.75e-19
C13374 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# -0.0489f
C13375 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__conb_1_51/HI 0.00675f
C13376 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__inv_1_54/Y 0.00498f
C13377 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_1_60/Y 1.33e-19
C13378 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00238f
C13379 sky130_fd_sc_hd__dfbbn_1_25/a_1672_329# V_GND 1.06e-19
C13380 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# sky130_fd_sc_hd__inv_1_11/Y 3.1e-21
C13381 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__inv_1_22/Y 0.0909f
C13382 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# -0.0178f
C13383 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_647_21# -0.00239f
C13384 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__inv_1_54/Y 1.47e-21
C13385 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__inv_1_75/A 0.0089f
C13386 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/Q_N 7.91e-19
C13387 FALLING_COUNTER.COUNT_SUB_DFF15.Q V_LOW 1.28f
C13388 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# sky130_fd_sc_hd__inv_1_17/Y 0.00173f
C13389 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/Q_N 2.34e-19
C13390 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# V_LOW 5.39e-19
C13391 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 3.86e-21
C13392 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# -0.0201f
C13393 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# -0.0078f
C13394 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0455f
C13395 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 7.12e-19
C13396 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# -3.46e-20
C13397 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 1.42e-32
C13398 sky130_fd_sc_hd__inv_1_86/Y sky130_fd_sc_hd__inv_1_93/A 3.49e-21
C13399 sky130_fd_sc_hd__conb_1_3/HI Reset 1.08e-20
C13400 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 4.62e-19
C13401 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# V_LOW -0.00266f
C13402 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_30/a_557_413# 1.77e-19
C13403 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__conb_1_46/HI 3.47e-19
C13404 sky130_fd_sc_hd__dfbbn_1_23/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.00406f
C13405 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_7/LO 0.00478f
C13406 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__inv_1_54/Y 6.53e-19
C13407 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.0245f
C13408 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 1.19e-19
C13409 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 7.97e-21
C13410 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_13/Y 3.94e-21
C13411 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00136f
C13412 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__inv_1_90/Y 0.0245f
C13413 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__conb_1_25/HI 0.0177f
C13414 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0151f
C13415 sky130_fd_sc_hd__conb_1_5/HI V_LOW 0.0285f
C13416 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00419f
C13417 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_71/A 0.0254f
C13418 sky130_fd_sc_hd__dfbbn_1_27/a_891_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.0012f
C13419 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# V_GND 0.00153f
C13420 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.98e-19
C13421 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 5.6e-19
C13422 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_28/Q_N 4.98e-19
C13423 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# V_LOW 0.00832f
C13424 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -0.00226f
C13425 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_83/Y 0.0164f
C13426 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# V_LOW 0.00598f
C13427 RISING_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 5.37e-20
C13428 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0451f
C13429 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 6e-19
C13430 sky130_fd_sc_hd__dfbbn_1_19/a_581_47# V_GND 1.91e-19
C13431 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# -5.42e-19
C13432 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 9.02e-19
C13433 RISING_COUNTER.COUNT_SUB_DFF2.Q V_LOW 3.63f
C13434 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 0.00104f
C13435 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__inv_1_23/Y 4.05e-20
C13436 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# 1.18e-19
C13437 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# sky130_fd_sc_hd__conb_1_46/HI 0.00102f
C13438 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__inv_1_47/Y 8.92e-19
C13439 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 3.61e-19
C13440 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 5.83e-21
C13441 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 8.03e-22
C13442 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0316f
C13443 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 3.01e-20
C13444 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_0/a_941_21# -1.42e-32
C13445 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# -0.00117f
C13446 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_0/a_381_47# -0.00811f
C13447 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__nand2_8_3/Y 6.94e-19
C13448 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 7.72e-19
C13449 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 2.26e-19
C13450 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# sky130_fd_sc_hd__inv_1_19/Y 0.0102f
C13451 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 0.00113f
C13452 sky130_fd_sc_hd__conb_1_4/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0517f
C13453 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_1672_329# 4.07e-20
C13454 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# Reset 0.00331f
C13455 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 9.57e-21
C13456 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0144f
C13457 sky130_fd_sc_hd__conb_1_14/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00232f
C13458 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/Q_N 6.25e-20
C13459 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# V_GND 0.00963f
C13460 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__conb_1_20/LO 0.00115f
C13461 sky130_fd_sc_hd__inv_1_78/A V_LOW 0.0842f
C13462 sky130_fd_sc_hd__dfbbn_1_27/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.00583f
C13463 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# sky130_fd_sc_hd__inv_1_19/Y 5.17e-20
C13464 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0542f
C13465 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0479f
C13466 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__inv_1_57/Y 4.02e-20
C13467 sky130_fd_sc_hd__dfbbn_1_47/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0166f
C13468 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__conb_1_20/HI -0.00838f
C13469 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00342f
C13470 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00401f
C13471 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 7.45e-19
C13472 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 0.00149f
C13473 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.00149f
C13474 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00386f
C13475 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_381_47# -0.00171f
C13476 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_791_47# -0.0122f
C13477 sky130_fd_sc_hd__conb_1_2/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 2.82e-19
C13478 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# CLOCK_GEN.SR_Op.Q 7.16e-19
C13479 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# -3.46e-20
C13480 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__conb_1_2/HI 0.0157f
C13481 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__inv_1_59/Y 5.69e-20
C13482 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 3.18e-19
C13483 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_28/Y 0.0443f
C13484 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_32/A 1.73e-19
C13485 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__inv_1_20/Y 5.85e-22
C13486 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__inv_1_4/Y 2.09e-19
C13487 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_4/LO 1.33e-19
C13488 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00612f
C13489 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__conb_1_37/HI 2.52e-21
C13490 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.05e-19
C13491 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# sky130_fd_sc_hd__inv_1_60/Y 1.83e-20
C13492 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# 1.58e-19
C13493 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 9.25e-20
C13494 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__inv_1_55/Y 2.18e-19
C13495 sky130_fd_sc_hd__conb_1_24/HI V_GND 0.104f
C13496 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# V_LOW -0.311f
C13497 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.97e-21
C13498 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 9.18e-19
C13499 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00109f
C13500 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0227f
C13501 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_75/Y 0.00205f
C13502 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_13/Q_N -6.48e-19
C13503 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 0.00982f
C13504 sky130_fd_sc_hd__inv_1_93/Y sky130_fd_sc_hd__inv_1_94/A 0.00514f
C13505 sky130_fd_sc_hd__inv_1_61/Y V_GND 0.116f
C13506 sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__inv_1_97/Y 0.519f
C13507 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0485f
C13508 sky130_fd_sc_hd__conb_1_7/HI V_GND 0.0192f
C13509 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__conb_1_46/HI 3.81e-20
C13510 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0063f
C13511 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 6.49e-21
C13512 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__inv_1_5/Y 0.00126f
C13513 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 1.62e-20
C13514 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_16_1/Y 0.00143f
C13515 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.12e-20
C13516 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__conb_1_48/HI 8.16e-19
C13517 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_16/Y 3.89e-20
C13518 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_76/A 0.00199f
C13519 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.05e-19
C13520 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# sky130_fd_sc_hd__inv_1_9/Y 6.17e-19
C13521 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 2.1e-20
C13522 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00534f
C13523 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# V_GND -0.00911f
C13524 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.26e-19
C13525 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# V_GND 0.00133f
C13526 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF10.Q 3.53e-19
C13527 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 0.00105f
C13528 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# sky130_fd_sc_hd__inv_1_53/Y 5.68e-19
C13529 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.03f
C13530 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF12.Q 8.2e-20
C13531 FULL_COUNTER.COUNT_SUB_DFF14.Q V_LOW 0.835f
C13532 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0707f
C13533 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_92/Y 0.0013f
C13534 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_13/HI 0.45f
C13535 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__inv_1_106/Y 3.76e-20
C13536 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__nand2_1_4/a_113_47# 7.29e-19
C13537 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 6.72e-21
C13538 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_22/LO 0.0539f
C13539 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.8e-20
C13540 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 1.14e-21
C13541 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 1.92e-22
C13542 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 5.12e-20
C13543 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.31e-19
C13544 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_1/a_791_47# 4.46e-20
C13545 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 4.38e-21
C13546 sky130_fd_sc_hd__dfbbn_1_5/a_1363_47# sky130_fd_sc_hd__inv_16_2/Y 2.48e-19
C13547 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_1_105/Y 0.109f
C13548 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__conb_1_21/HI 0.0248f
C13549 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 5.13e-20
C13550 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.6e-21
C13551 sky130_fd_sc_hd__dfbbn_1_9/a_581_47# sky130_fd_sc_hd__inv_1_19/Y 1.39e-19
C13552 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# 3.59e-19
C13553 sky130_fd_sc_hd__dfbbn_1_31/Q_N Reset 0.0176f
C13554 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0856f
C13555 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__conb_1_5/HI 2.17e-20
C13556 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0059f
C13557 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# V_GND 0.00248f
C13558 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/Q_N -4.24e-20
C13559 sky130_fd_sc_hd__dfbbn_1_8/Q_N sky130_fd_sc_hd__inv_1_19/Y 5.39e-21
C13560 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__conb_1_28/HI 4.73e-19
C13561 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__conb_1_20/HI -1.1e-19
C13562 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.16f
C13563 RISING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_59/Y 2.07e-20
C13564 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# -1.44e-20
C13565 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# CLOCK_GEN.SR_Op.Q 4.32e-22
C13566 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__conb_1_44/HI 3.48e-19
C13567 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 7.27e-20
C13568 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0.0123f
C13569 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 6.69e-21
C13570 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__inv_1_58/Y 1.46e-19
C13571 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__conb_1_23/HI -0.0014f
C13572 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.0919f
C13573 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 3.93e-19
C13574 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__inv_1_55/Y 3.67e-19
C13575 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 3.43e-20
C13576 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 3.98e-19
C13577 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 1.35e-19
C13578 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# sky130_fd_sc_hd__inv_1_53/Y 0.0179f
C13579 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 1.65e-20
C13580 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__nand2_8_9/Y 1.83e-20
C13581 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__conb_1_25/HI 0.0245f
C13582 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.0132f
C13583 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.026f
C13584 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 6.84e-20
C13585 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 9.29e-20
C13586 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# 9.98e-19
C13587 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF8.Q 0.196f
C13588 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.4e-19
C13589 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_101/Y 0.111f
C13590 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 7.36e-19
C13591 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_20/LO 1.06e-19
C13592 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 7.29e-20
C13593 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0137f
C13594 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.6e-19
C13595 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 2.28e-21
C13596 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.27e-19
C13597 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# CLOCK_GEN.SR_Op.Q 0.0139f
C13598 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# V_LOW -0.00389f
C13599 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__inv_1_11/Y 1.26e-19
C13600 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0239f
C13601 sky130_fd_sc_hd__dfbbn_1_21/Q_N RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00255f
C13602 sky130_fd_sc_hd__dfbbn_1_39/a_1672_329# V_GND 2.44e-19
C13603 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_1_105/Y 0.0256f
C13604 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# sky130_fd_sc_hd__inv_1_54/Y 0.00651f
C13605 sky130_fd_sc_hd__conb_1_28/LO sky130_fd_sc_hd__inv_16_1/Y 1.13e-20
C13606 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 5.04e-21
C13607 sky130_fd_sc_hd__dfbbn_1_30/Q_N V_GND -0.00201f
C13608 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 8.79e-21
C13609 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 6.25e-19
C13610 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0.00449f
C13611 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 4.81e-21
C13612 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/Q_N -4.33e-20
C13613 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 2.39e-20
C13614 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.46e-20
C13615 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 4.62e-19
C13616 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 3.16e-19
C13617 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.0197f
C13618 FALLING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_103/Y 8.81e-20
C13619 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# sky130_fd_sc_hd__inv_1_18/Y 0.00326f
C13620 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 5.17e-19
C13621 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# V_GND 9.21e-19
C13622 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# sky130_fd_sc_hd__conb_1_6/HI 7.99e-20
C13623 sky130_fd_sc_hd__conb_1_39/LO sky130_fd_sc_hd__inv_16_1/Y 7.46e-19
C13624 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/Q_N -9.56e-20
C13625 sky130_fd_sc_hd__inv_1_95/Y V_LOW 0.158f
C13626 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 7.33e-21
C13627 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0151f
C13628 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__conb_1_22/HI 1.12e-20
C13629 sky130_fd_sc_hd__dfbbn_1_21/Q_N sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.69e-20
C13630 sky130_fd_sc_hd__dfbbn_1_16/a_581_47# sky130_fd_sc_hd__conb_1_5/HI 7.95e-20
C13631 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0367f
C13632 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 0.00633f
C13633 sky130_fd_sc_hd__dfbbn_1_35/Q_N V_GND 0.00168f
C13634 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0292f
C13635 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.00155f
C13636 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__conb_1_21/HI 3.53e-20
C13637 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__conb_1_20/HI -1.59e-19
C13638 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# sky130_fd_sc_hd__inv_1_8/Y 7.55e-20
C13639 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 0.00202f
C13640 sky130_fd_sc_hd__dfbbn_1_38/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.00717f
C13641 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 5.83e-20
C13642 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0.0013f
C13643 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__conb_1_4/HI 0.0134f
C13644 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_1/a_113_47# 5.21e-19
C13645 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0056f
C13646 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_50/a_27_47# 2.13e-20
C13647 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# -0.00458f
C13648 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# -0.0106f
C13649 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_41/a_381_47# -3.04e-19
C13650 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# -6.23e-21
C13651 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 1.01e-20
C13652 FULL_COUNTER.COUNT_SUB_DFF0.Q Reset 6.16e-19
C13653 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_39/LO 2.87e-20
C13654 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_42/LO 0.0462f
C13655 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0127f
C13656 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_18/HI 1.18e-19
C13657 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_1_98/Y 1.72e-19
C13658 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# V_GND 0.0617f
C13659 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 2.65e-20
C13660 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 5.05e-19
C13661 sky130_fd_sc_hd__inv_1_81/Y Reset 0.0319f
C13662 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__conb_1_18/HI -0.00108f
C13663 FALLING_COUNTER.COUNT_SUB_DFF7.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 4.84e-21
C13664 sky130_fd_sc_hd__inv_1_92/Y sky130_fd_sc_hd__inv_1_86/Y 0.00527f
C13665 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__conb_1_23/HI -0.0127f
C13666 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 3.89e-20
C13667 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 0.0123f
C13668 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__conb_1_41/HI 4.71e-20
C13669 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# sky130_fd_sc_hd__conb_1_25/HI -0.0125f
C13670 sky130_fd_sc_hd__dfbbn_1_28/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.00278f
C13671 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_16_2/Y 0.0541f
C13672 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.5e-19
C13673 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_75/Y 1.23e-20
C13674 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_7/Y 1.08e-20
C13675 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 0.0245f
C13676 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__nand3_1_2/B 6.72e-20
C13677 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__conb_1_30/HI -0.0155f
C13678 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_381_47# -2.53e-20
C13679 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 6.84e-21
C13680 sky130_fd_sc_hd__inv_16_1/Y sky130_fd_sc_hd__inv_1_108/Y 0.103f
C13681 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_74/Y 9.88e-19
C13682 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__conb_1_11/HI 5.54e-21
C13683 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 0.578f
C13684 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__conb_1_24/HI 0.00126f
C13685 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 9.82e-21
C13686 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 3.2e-21
C13687 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 5.1e-21
C13688 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 1.53e-20
C13689 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__conb_1_18/HI 8.83e-19
C13690 sky130_fd_sc_hd__conb_1_37/HI V_GND 0.286f
C13691 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__conb_1_22/HI 0.00402f
C13692 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 7.61e-20
C13693 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_4/LO 3.38e-20
C13694 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_11/LO 0.0238f
C13695 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00464f
C13696 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_1_105/Y 0.0194f
C13697 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.34e-20
C13698 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__inv_1_76/A 0.00758f
C13699 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_93/A 0.292f
C13700 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_41/a_27_47# 2.32e-19
C13701 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_16/HI -7.53e-19
C13702 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__conb_1_39/HI 5.84e-21
C13703 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__inv_1_9/Y 6.7e-21
C13704 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 2.69e-19
C13705 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 3.16e-19
C13706 sky130_fd_sc_hd__inv_1_17/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0252f
C13707 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__nand2_8_9/Y 3.52e-20
C13708 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# V_LOW 1.38e-19
C13709 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00492f
C13710 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# V_LOW 0.0204f
C13711 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_193_47# 0.00196f
C13712 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 0.00173f
C13713 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 7.59e-21
C13714 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# sky130_fd_sc_hd__inv_16_0/Y 3.94e-19
C13715 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 6.86e-20
C13716 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.03e-19
C13717 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# V_LOW -0.00554f
C13718 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00436f
C13719 sky130_fd_sc_hd__dfbbn_1_8/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00113f
C13720 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.38e-19
C13721 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# -6.22e-19
C13722 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# -0.00464f
C13723 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# -6.23e-21
C13724 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.063f
C13725 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0197f
C13726 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0218f
C13727 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_891_329# 9.3e-19
C13728 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00202f
C13729 sky130_fd_sc_hd__nand2_8_8/a_27_47# CLOCK_GEN.SR_Op.Q 0.0379f
C13730 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 0.00407f
C13731 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 3.81e-19
C13732 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_50/A 0.0207f
C13733 sky130_fd_sc_hd__inv_1_66/Y sky130_fd_sc_hd__inv_1_93/A 0.00159f
C13734 sky130_fd_sc_hd__dfbbn_1_2/a_557_413# V_LOW 3.56e-20
C13735 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__inv_1_57/Y 0.00796f
C13736 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# 8.88e-20
C13737 sky130_fd_sc_hd__dfbbn_1_37/a_1112_329# V_GND 0.00104f
C13738 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.104f
C13739 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 7.64e-19
C13740 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__inv_1_99/Y 0.00113f
C13741 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# V_GND 0.00589f
C13742 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# V_LOW 0.00684f
C13743 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0137f
C13744 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__conb_1_46/LO 8.84e-20
C13745 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0218f
C13746 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__inv_1_76/A 4.43e-19
C13747 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# V_LOW 0.0131f
C13748 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# V_GND 0.00372f
C13749 sky130_fd_sc_hd__inv_1_93/A V_GND 0.439f
C13750 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# sky130_fd_sc_hd__conb_1_21/HI -2.6e-20
C13751 sky130_fd_sc_hd__conb_1_26/LO V_LOW 0.143f
C13752 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__conb_1_40/HI 0.00621f
C13753 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 5.82e-20
C13754 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__conb_1_35/HI 0.415f
C13755 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 7.14e-20
C13756 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 4.49e-19
C13757 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 1.46e-19
C13758 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 5.31e-19
C13759 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 5.13e-19
C13760 FULL_COUNTER.COUNT_SUB_DFF1.Q V_LOW 2.16f
C13761 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_9/HI 0.00539f
C13762 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 6.39e-19
C13763 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# sky130_fd_sc_hd__inv_1_6/Y 3.75e-21
C13764 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_1_107/Y 0.00345f
C13765 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_13/HI 7.82e-21
C13766 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__nand2_8_2/A 0.00849f
C13767 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 9.87e-19
C13768 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_16_2/Y 0.0661f
C13769 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 5.55e-19
C13770 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__inv_1_98/Y 9.37e-21
C13771 sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# V_GND 1.99e-19
C13772 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# sky130_fd_sc_hd__conb_1_18/HI -4.01e-20
C13773 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# V_GND 5.15e-19
C13774 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.48e-19
C13775 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__conb_1_38/HI 0.0284f
C13776 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# V_LOW 0.00649f
C13777 sky130_fd_sc_hd__dfbbn_1_50/a_891_329# V_GND 4.5e-19
C13778 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.9e-19
C13779 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 2.62e-19
C13780 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0102f
C13781 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# V_LOW 2.64e-19
C13782 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_23/HI 0.0113f
C13783 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_1_98/Y 2.23e-19
C13784 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF1.Q 0.187f
C13785 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_71/Y 0.00904f
C13786 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0102f
C13787 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# sky130_fd_sc_hd__inv_1_106/Y 7.97e-21
C13788 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_22/a_381_47# -3.79e-20
C13789 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_22/a_1112_329# -4.66e-20
C13790 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# -0.00117f
C13791 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# -0.00367f
C13792 sky130_fd_sc_hd__inv_1_32/Y V_GND 0.0853f
C13793 RISING_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 5.36e-21
C13794 sky130_fd_sc_hd__inv_1_46/Y V_GND 0.121f
C13795 FALLING_COUNTER.COUNT_SUB_DFF14.Q V_LOW 1.72f
C13796 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 2.41e-20
C13797 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 4.06e-19
C13798 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.32e-21
C13799 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# sky130_fd_sc_hd__conb_1_30/HI -9.57e-19
C13800 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# -1.44e-20
C13801 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 9.35e-21
C13802 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__conb_1_26/HI 1.86e-19
C13803 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# -6.23e-21
C13804 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__dfbbn_1_31/a_941_21# -9.88e-20
C13805 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_31/a_381_47# -0.00464f
C13806 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# V_LOW 7.94e-19
C13807 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 3.67e-22
C13808 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# V_GND -0.00496f
C13809 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_67/Y 0.0225f
C13810 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# sky130_fd_sc_hd__conb_1_22/HI 0.00217f
C13811 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__conb_1_44/HI 0.00257f
C13812 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF6.Q 4.06e-21
C13813 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# V_GND -0.00443f
C13814 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_1112_329# -0.00336f
C13815 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_381_47# -3.79e-20
C13816 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF14.Q 2.42e-19
C13817 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_41/a_1340_413# 1.01e-20
C13818 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# sky130_fd_sc_hd__conb_1_16/HI 0.00624f
C13819 sky130_fd_sc_hd__inv_1_10/Y V_GND 0.0982f
C13820 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# sky130_fd_sc_hd__inv_1_9/Y 3.16e-19
C13821 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 4.28e-20
C13822 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0.00616f
C13823 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00131f
C13824 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_72/Y 0.0156f
C13825 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0.0151f
C13826 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_40/HI 0.0356f
C13827 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 8.29e-20
C13828 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 5.67e-19
C13829 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 4.06e-21
C13830 sky130_fd_sc_hd__conb_1_2/LO FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0113f
C13831 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.36e-20
C13832 sky130_fd_sc_hd__dfbbn_1_0/a_557_413# V_GND 1.83e-19
C13833 sky130_fd_sc_hd__inv_1_93/A sky130_fd_sc_hd__nand3_1_1/Y 8.28e-19
C13834 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_63/Y 1.53e-20
C13835 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.58e-19
C13836 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_6/HI 5.24e-19
C13837 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__conb_1_39/HI 1.85e-19
C13838 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0558f
C13839 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00106f
C13840 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF0.Q 5.3e-21
C13841 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00525f
C13842 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 4.45e-19
C13843 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.0014f
C13844 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# sky130_fd_sc_hd__inv_1_18/Y 0.00233f
C13845 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00339f
C13846 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_891_329# 2.24e-19
C13847 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_1112_329# -4.66e-20
C13848 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__conb_1_18/HI 6.71e-20
C13849 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/Q_N 5.7e-19
C13850 sky130_fd_sc_hd__nand3_1_1/a_193_47# V_GND 3.27e-19
C13851 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__inv_1_99/Y 8.44e-19
C13852 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# V_GND 2.65e-19
C13853 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# -7.77e-19
C13854 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -0.00556f
C13855 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF0.Q 2.67e-20
C13856 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00818f
C13857 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# V_LOW 4.14e-20
C13858 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00185f
C13859 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_32/HI 0.0277f
C13860 sky130_fd_sc_hd__dfbbn_1_33/a_891_329# sky130_fd_sc_hd__conb_1_35/HI 8.25e-19
C13861 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# V_LOW 4.7e-20
C13862 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# V_GND 0.00212f
C13863 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__inv_1_54/Y 4.43e-21
C13864 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 1.28e-20
C13865 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# -3.06e-20
C13866 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# -0.00631f
C13867 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# Reset 5.59e-19
C13868 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__inv_1_23/Y 0.0047f
C13869 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 8.27e-19
C13870 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 1.25e-20
C13871 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__inv_1_47/Y 4.56e-21
C13872 sky130_fd_sc_hd__dfbbn_1_51/a_1159_47# sky130_fd_sc_hd__conb_1_40/HI 2.09e-19
C13873 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 4.01e-20
C13874 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/Q_N 0.0014f
C13875 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_27/LO 0.0537f
C13876 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 5.19e-21
C13877 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 6.01e-21
C13878 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/Q_N -7.69e-20
C13879 sky130_fd_sc_hd__inv_1_72/A V_LOW 0.248f
C13880 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0127f
C13881 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__inv_1_107/Y 0.0295f
C13882 FULL_COUNTER.COUNT_SUB_DFF15.Q V_GND 1.02f
C13883 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00337f
C13884 sky130_fd_sc_hd__conb_1_6/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 2.19e-21
C13885 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.01f
C13886 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_102/Y 0.0352f
C13887 RISING_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 7.61e-20
C13888 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 1.46f
C13889 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 3.64e-19
C13890 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__conb_1_38/HI -0.0121f
C13891 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_85/Y 7.76e-20
C13892 sky130_fd_sc_hd__dfbbn_1_45/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.37e-19
C13893 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_96/Y 2.62e-19
C13894 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.00257f
C13895 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__inv_1_98/Y 0.0017f
C13896 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.4e-20
C13897 sky130_fd_sc_hd__dfbbn_1_20/a_891_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00162f
C13898 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.1e-20
C13899 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/Q_N 0.0114f
C13900 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 5.1e-21
C13901 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_94/A 4.76e-19
C13902 sky130_fd_sc_hd__dfbbn_1_26/Q_N sky130_fd_sc_hd__conb_1_30/HI -1.85e-19
C13903 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 1.94e-21
C13904 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__conb_1_47/HI 6.02e-20
C13905 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# -2.52e-19
C13906 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -0.0116f
C13907 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__conb_1_17/HI 2.52e-19
C13908 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# V_LOW 0.0101f
C13909 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00146f
C13910 sky130_fd_sc_hd__conb_1_28/LO V_LOW 0.0988f
C13911 sky130_fd_sc_hd__conb_1_4/HI V_LOW 0.186f
C13912 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.24e-21
C13913 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# V_GND -0.00504f
C13914 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_16_1/Y 2.18e-20
C13915 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00505f
C13916 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# V_GND -0.00515f
C13917 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_31/Y 0.156f
C13918 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__inv_1_55/Y 0.00443f
C13919 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# V_LOW -0.0042f
C13920 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0.00217f
C13921 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# V_LOW 0.0168f
C13922 sky130_fd_sc_hd__dfbbn_1_10/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00288f
C13923 sky130_fd_sc_hd__conb_1_39/LO V_LOW 0.0993f
C13924 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# -4.66e-20
C13925 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# -3.79e-20
C13926 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# sky130_fd_sc_hd__conb_1_40/HI 0.00758f
C13927 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__inv_1_66/Y 0.00937f
C13928 sky130_fd_sc_hd__nand3_1_1/a_193_47# sky130_fd_sc_hd__nand3_1_1/Y 6.73e-19
C13929 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__conb_1_29/LO 0.00107f
C13930 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0252f
C13931 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.33f
C13932 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_30/LO 0.00114f
C13933 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_34/a_941_21# 5.93e-20
C13934 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0476f
C13935 sky130_fd_sc_hd__dfbbn_1_25/a_557_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 4.31e-19
C13936 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF0.Q 6.71e-21
C13937 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 7.99e-19
C13938 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# sky130_fd_sc_hd__conb_1_39/HI -5.61e-19
C13939 sky130_fd_sc_hd__dfbbn_1_20/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 3.35e-19
C13940 sky130_fd_sc_hd__dfbbn_1_50/Q_N FALLING_COUNTER.COUNT_SUB_DFF0.Q 8.5e-19
C13941 sky130_fd_sc_hd__inv_1_78/A sky130_fd_sc_hd__inv_1_80/A 0.00409f
C13942 sky130_fd_sc_hd__inv_1_94/A V_GND 0.718f
C13943 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 4.35e-20
C13944 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__conb_1_26/HI 1.14e-20
C13945 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0144f
C13946 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.06e-20
C13947 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_1_100/Y 2.8e-20
C13948 sky130_fd_sc_hd__dfbbn_1_12/a_581_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.35e-20
C13949 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 0.0295f
C13950 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# V_GND 0.00158f
C13951 sky130_fd_sc_hd__dfbbn_1_41/a_557_413# V_GND 2.71e-19
C13952 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# FULL_COUNTER.COUNT_SUB_DFF15.Q 4.57e-19
C13953 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# -1.66e-19
C13954 sky130_fd_sc_hd__inv_1_19/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 9.03e-20
C13955 sky130_fd_sc_hd__dfbbn_1_38/Q_N V_LOW 5.07e-19
C13956 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__conb_1_32/HI -0.0122f
C13957 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# V_LOW 0.0274f
C13958 sky130_fd_sc_hd__dfbbn_1_23/Q_N V_GND 0.00142f
C13959 sky130_fd_sc_hd__dfbbn_1_50/Q_N V_LOW -0.00509f
C13960 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__inv_1_112/Y 4.51e-19
C13961 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0396f
C13962 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 7.69e-21
C13963 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__nand3_1_2/Y 0.285f
C13964 sky130_fd_sc_hd__conb_1_0/HI sky130_fd_sc_hd__conb_1_2/HI 0.00427f
C13965 sky130_fd_sc_hd__conb_1_35/LO sky130_fd_sc_hd__conb_1_37/HI 8.84e-20
C13966 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__nand2_8_2/A 6.85e-20
C13967 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00697f
C13968 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_381_47# -0.00441f
C13969 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_1_11/Y 6.37e-19
C13970 sky130_fd_sc_hd__conb_1_2/LO sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 1.05e-19
C13971 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# Reset 0.00233f
C13972 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 8.48e-21
C13973 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__nand2_8_3/Y 8.58e-20
C13974 sky130_fd_sc_hd__dfbbn_1_24/a_557_413# V_GND 2.12e-19
C13975 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.47e-19
C13976 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__conb_1_11/HI 2.27e-20
C13977 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__inv_1_103/Y 1.99e-21
C13978 RISING_COUNTER.COUNT_SUB_DFF0.Q Reset 0.0271f
C13979 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__inv_1_98/Y 0.00575f
C13980 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.43e-21
C13981 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 5.88e-20
C13982 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_2/a_193_47# 1.97e-35
C13983 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/Q_N -7.69e-20
C13984 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_473_413# -0.0222f
C13985 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -0.00369f
C13986 sky130_fd_sc_hd__inv_1_108/Y V_LOW 0.0554f
C13987 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 2.31e-20
C13988 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.83e-20
C13989 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# CLOCK_GEN.SR_Op.Q 8.03e-20
C13990 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__conb_1_47/HI 2.86e-20
C13991 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0115f
C13992 sky130_fd_sc_hd__inv_1_59/Y sky130_fd_sc_hd__inv_1_60/Y 0.00372f
C13993 transmission_gate_0/GN V_GND 0.00264f
C13994 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00107f
C13995 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# -1.76e-19
C13996 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# -7.17e-20
C13997 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_92/Y 8.02e-20
C13998 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# sky130_fd_sc_hd__conb_1_17/HI 2.43e-19
C13999 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00106f
C14000 sky130_fd_sc_hd__dfbbn_1_27/Q_N V_GND -0.00767f
C14001 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF13.Q 3.49e-21
C14002 sky130_fd_sc_hd__dfbbn_1_47/Q_N V_GND -0.00767f
C14003 sky130_fd_sc_hd__conb_1_36/LO sky130_fd_sc_hd__inv_1_108/Y 2.42e-19
C14004 RISING_COUNTER.COUNT_SUB_DFF9.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.903f
C14005 sky130_fd_sc_hd__inv_1_94/A sky130_fd_sc_hd__nand3_1_1/Y 0.0178f
C14006 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# -3.04e-19
C14007 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# -0.00133f
C14008 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# V_LOW -4.72e-19
C14009 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.21e-20
C14010 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# V_LOW -0.00136f
C14011 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 1.52e-19
C14012 sky130_fd_sc_hd__dfbbn_1_47/a_1112_329# sky130_fd_sc_hd__inv_1_57/Y 0.00179f
C14013 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 3.13e-21
C14014 sky130_fd_sc_hd__dfbbn_1_17/Q_N FULL_COUNTER.COUNT_SUB_DFF8.Q 1.9e-20
C14015 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 6.05e-20
C14016 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.28e-20
C14017 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__conb_1_42/LO 8.84e-20
C14018 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__conb_1_24/LO 2.83e-21
C14019 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0.00599f
C14020 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0.00132f
C14021 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0.00142f
C14022 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 0.00105f
C14023 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__inv_1_102/Y 2.1e-21
C14024 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 0.00725f
C14025 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_1_5/Y 1.15e-19
C14026 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# V_LOW -0.0633f
C14027 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 7.62e-20
C14028 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 0.00542f
C14029 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__conb_1_26/HI 5.52e-20
C14030 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.97e-19
C14031 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__conb_1_4/HI 0.0174f
C14032 sky130_fd_sc_hd__inv_1_92/Y V_GND 0.563f
C14033 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 2.86e-19
C14034 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 1.62e-19
C14035 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 2.27e-19
C14036 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 7.9e-19
C14037 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# V_GND 0.00836f
C14038 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# V_GND 0.00122f
C14039 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 1.86e-20
C14040 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0315f
C14041 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# V_LOW 0.00789f
C14042 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_105/Y 0.0368f
C14043 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_32/HI 4.56e-21
C14044 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_891_329# 1.48e-20
C14045 RISING_COUNTER.COUNT_SUB_DFF2.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00113f
C14046 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_17/HI 9.92e-19
C14047 sky130_fd_sc_hd__dfbbn_1_9/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00461f
C14048 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# sky130_fd_sc_hd__inv_1_107/Y 9.54e-19
C14049 sky130_fd_sc_hd__conb_1_1/LO V_LOW 0.0977f
C14050 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.95e-22
C14051 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_31/HI 0.35f
C14052 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_57/Y 4.98e-21
C14053 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# V_GND -5.48e-19
C14054 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__conb_1_0/HI 1.09e-19
C14055 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__conb_1_1/HI 0.0114f
C14056 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 5.51e-20
C14057 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# V_GND -0.00547f
C14058 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.72e-20
C14059 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# sky130_fd_sc_hd__inv_1_103/Y 2.5e-20
C14060 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__conb_1_36/HI 0.00179f
C14061 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# -1.44e-20
C14062 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# Reset 4.28e-19
C14063 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.053f
C14064 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_581_47# 1.06e-19
C14065 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# sky130_fd_sc_hd__inv_1_61/Y 0.00983f
C14066 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 9.9e-19
C14067 sky130_fd_sc_hd__inv_16_0/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 0.178f
C14068 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_57/Y 0.00261f
C14069 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__inv_1_63/Y 2.31e-20
C14070 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# sky130_fd_sc_hd__conb_1_34/HI 0.00134f
C14071 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.95e-20
C14072 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0139f
C14073 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__conb_1_42/HI 0.0213f
C14074 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.06e-20
C14075 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_45/HI 2.87e-19
C14076 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__conb_1_38/HI 1.03e-19
C14077 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.19e-20
C14078 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__inv_1_59/Y 8.57e-19
C14079 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# sky130_fd_sc_hd__conb_1_24/HI -0.0757f
C14080 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_2/a_791_47# 5.78e-20
C14081 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0.0326f
C14082 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0125f
C14083 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 2.12e-19
C14084 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 0.0138f
C14085 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__conb_1_2/HI 0.00138f
C14086 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# -0.0103f
C14087 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# -0.00251f
C14088 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__inv_1_102/Y 3.49e-19
C14089 sky130_fd_sc_hd__dfbbn_1_12/Q_N sky130_fd_sc_hd__conb_1_17/HI 4.38e-20
C14090 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 4.02e-19
C14091 FULL_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_6/HI 0.044f
C14092 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 1.29e-19
C14093 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_108/Y 1.3e-19
C14094 sky130_fd_sc_hd__inv_1_48/Y V_GND 0.0264f
C14095 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 1.53e-20
C14096 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_1_4/Y 1.72e-20
C14097 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_102/Y 2.93e-20
C14098 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 6.09e-20
C14099 sky130_fd_sc_hd__inv_1_71/A Reset 0.0252f
C14100 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 1.03e-21
C14101 sky130_fd_sc_hd__dfbbn_1_48/a_557_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00133f
C14102 sky130_fd_sc_hd__inv_1_95/Y sky130_fd_sc_hd__inv_1_80/A 1.07e-20
C14103 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 2.62e-20
C14104 FULL_COUNTER.COUNT_SUB_DFF2.Q V_LOW 0.786f
C14105 sky130_fd_sc_hd__conb_1_10/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 9.87e-21
C14106 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 0.0278f
C14107 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__conb_1_13/HI 1.72e-20
C14108 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.49e-20
C14109 sky130_fd_sc_hd__dfbbn_1_45/Q_N FALLING_COUNTER.COUNT_SUB_DFF8.Q 4.27e-19
C14110 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_13/Y 5.41e-22
C14111 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 5.85e-20
C14112 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# V_LOW -0.00121f
C14113 sky130_fd_sc_hd__inv_1_111/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0725f
C14114 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_1340_413# 8.48e-19
C14115 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_581_47# 5.8e-19
C14116 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# V_LOW -2.68e-19
C14117 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 3.82e-19
C14118 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__conb_1_26/HI 4.76e-20
C14119 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_42/HI 0.0181f
C14120 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 1.54e-22
C14121 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# V_GND 0.00382f
C14122 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_791_47# 2.75e-20
C14123 sky130_fd_sc_hd__dfbbn_1_33/Q_N V_GND -0.00224f
C14124 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0399f
C14125 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__inv_1_58/Y 5.15e-19
C14126 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 4.37e-20
C14127 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__conb_1_38/HI 4.77e-19
C14128 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_473_413# 0.00109f
C14129 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# sky130_fd_sc_hd__inv_1_107/Y 1.85e-19
C14130 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0463f
C14131 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.002f
C14132 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__conb_1_10/HI -0.00143f
C14133 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 0.00267f
C14134 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_39/A 0.652f
C14135 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0238f
C14136 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_891_329# 7.79e-19
C14137 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# V_LOW -0.0213f
C14138 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# V_GND -0.00483f
C14139 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_473_413# -3.86e-20
C14140 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# -0.00408f
C14141 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__conb_1_10/HI 8.86e-20
C14142 sky130_fd_sc_hd__dfbbn_1_39/Q_N FALLING_COUNTER.COUNT_SUB_DFF11.Q 9.66e-20
C14143 sky130_fd_sc_hd__dfbbn_1_3/a_1363_47# sky130_fd_sc_hd__conb_1_0/HI -2.6e-20
C14144 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# sky130_fd_sc_hd__conb_1_36/HI -2.1e-20
C14145 sky130_fd_sc_hd__dfbbn_1_32/a_1363_47# V_GND -3.83e-19
C14146 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 3.65e-20
C14147 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# sky130_fd_sc_hd__inv_1_103/Y 2.66e-21
C14148 sky130_fd_sc_hd__dfbbn_1_40/a_1159_47# sky130_fd_sc_hd__conb_1_36/HI 0.00152f
C14149 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__conb_1_25/LO 8.84e-20
C14150 sky130_fd_sc_hd__dfbbn_1_39/a_1159_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 5.18e-19
C14151 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 0.00808f
C14152 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.213f
C14153 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# sky130_fd_sc_hd__conb_1_51/HI 7.77e-19
C14154 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__conb_1_48/LO 8.81e-20
C14155 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# sky130_fd_sc_hd__conb_1_11/HI 0.00519f
C14156 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# V_LOW 0.0325f
C14157 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__conb_1_6/LO 2.53e-20
C14158 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# V_GND 0.0215f
C14159 sky130_fd_sc_hd__conb_1_37/LO FALLING_COUNTER.COUNT_SUB_DFF8.Q 3.8e-19
C14160 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# sky130_fd_sc_hd__conb_1_42/HI 0.00516f
C14161 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# sky130_fd_sc_hd__conb_1_45/HI 1.3e-19
C14162 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 0.00607f
C14163 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.11e-19
C14164 sky130_fd_sc_hd__dfbbn_1_43/a_1672_329# sky130_fd_sc_hd__inv_1_59/Y 7.32e-19
C14165 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# sky130_fd_sc_hd__inv_1_10/Y 0.00525f
C14166 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# V_GND -0.00441f
C14167 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__conb_1_40/HI 5.02e-19
C14168 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.0055f
C14169 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.96e-19
C14170 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 6.09e-21
C14171 sky130_fd_sc_hd__dfbbn_1_46/a_581_47# sky130_fd_sc_hd__inv_16_1/Y 0.00181f
C14172 sky130_fd_sc_hd__conb_1_29/HI V_LOW 0.014f
C14173 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# -9.41e-19
C14174 sky130_fd_sc_hd__dfbbn_1_30/a_581_47# sky130_fd_sc_hd__inv_1_102/Y 2.34e-19
C14175 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_581_47# 1.69e-19
C14176 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.47e-20
C14177 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 9.61e-22
C14178 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.44e-20
C14179 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# V_GND 0.00948f
C14180 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 3.5e-21
C14181 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# V_GND 0.0556f
C14182 FULL_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_12/HI 5.67e-20
C14183 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# sky130_fd_sc_hd__inv_1_108/Y 2.06e-19
C14184 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00541f
C14185 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# V_GND 2.89e-19
C14186 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# sky130_fd_sc_hd__inv_1_21/Y 0.00113f
C14187 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__inv_1_15/Y 9.96e-20
C14188 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/Q_N -9.56e-20
C14189 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 0.00697f
C14190 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# V_LOW 0.0243f
C14191 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 7.39e-21
C14192 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0698f
C14193 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0332f
C14194 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 9.59e-19
C14195 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# -1.03e-19
C14196 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_473_413# -3.86e-20
C14197 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.15e-20
C14198 FALLING_COUNTER.COUNT_SUB_DFF6.Q Reset 0.00689f
C14199 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_70/Y 0.00144f
C14200 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 8.8e-21
C14201 sky130_fd_sc_hd__inv_1_32/A V_SENSE 0.0961f
C14202 sky130_fd_sc_hd__conb_1_19/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 1.48e-20
C14203 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.59e-21
C14204 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 9.75e-19
C14205 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 1.68e-19
C14206 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 2.52e-19
C14207 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__conb_1_22/HI 6.64e-19
C14208 sky130_fd_sc_hd__dfbbn_1_2/Q_N sky130_fd_sc_hd__conb_1_2/HI 0.00162f
C14209 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__conb_1_42/HI -0.0122f
C14210 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__inv_1_98/Y 1.16e-22
C14211 sky130_fd_sc_hd__conb_1_3/LO CLOCK_GEN.SR_Op.Q 1.56e-20
C14212 sky130_fd_sc_hd__dfbbn_1_28/Q_N V_GND 0.00296f
C14213 sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00708f
C14214 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# V_GND -0.00527f
C14215 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_381_47# -0.00516f
C14216 sky130_fd_sc_hd__dfbbn_1_27/Q_N RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0154f
C14217 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__inv_1_22/Y 0.018f
C14218 sky130_fd_sc_hd__conb_1_49/HI FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00389f
C14219 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 1.77e-19
C14220 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 7.02e-19
C14221 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# V_LOW 2.26e-20
C14222 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.95e-20
C14223 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# V_LOW 0.00828f
C14224 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__conb_1_27/HI 0.0232f
C14225 sky130_fd_sc_hd__inv_1_21/Y V_LOW 0.245f
C14226 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1159_47# 0.00105f
C14227 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0131f
C14228 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 0.00105f
C14229 sky130_fd_sc_hd__conb_1_27/LO CLOCK_GEN.SR_Op.Q 2.47e-19
C14230 sky130_fd_sc_hd__dfbbn_1_6/a_1159_47# sky130_fd_sc_hd__conb_1_10/HI -9.78e-19
C14231 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__inv_1_60/Y 8.14e-19
C14232 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# V_LOW -0.0203f
C14233 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00268f
C14234 sky130_fd_sc_hd__conb_1_18/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 7.63e-19
C14235 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# V_LOW -1.01e-19
C14236 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_56/Y 1.82e-21
C14237 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_1340_413# -9.41e-19
C14238 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# sky130_fd_sc_hd__conb_1_36/HI -0.01f
C14239 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 0.0102f
C14240 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# V_LOW -4e-20
C14241 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__conb_1_47/HI 8.16e-19
C14242 sky130_fd_sc_hd__dfbbn_1_11/a_1112_329# sky130_fd_sc_hd__inv_1_22/Y 5.15e-21
C14243 sky130_fd_sc_hd__inv_1_70/A sky130_fd_sc_hd__nand2_8_9/Y 0.00331f
C14244 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.61e-19
C14245 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 0.00268f
C14246 sky130_fd_sc_hd__conb_1_20/LO V_GND 0.00105f
C14247 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 3.89e-19
C14248 sky130_fd_sc_hd__dfbbn_1_29/a_1340_413# V_LOW 2.94e-20
C14249 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# V_GND 0.00202f
C14250 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# V_GND 0.00106f
C14251 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_381_47# -2.53e-20
C14252 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# V_LOW -9.15e-19
C14253 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# V_LOW 4.8e-20
C14254 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# -0.00539f
C14255 sky130_fd_sc_hd__dfbbn_1_12/a_557_413# V_GND 1.76e-19
C14256 sky130_fd_sc_hd__inv_1_13/Y FULL_COUNTER.COUNT_SUB_DFF5.Q 0.172f
C14257 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 9.92e-20
C14258 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_76/A 0.00506f
C14259 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 4.73e-19
C14260 sky130_fd_sc_hd__inv_1_69/Y sky130_fd_sc_hd__inv_1_68/Y 0.00125f
C14261 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# V_GND -0.00162f
C14262 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# -5.54e-21
C14263 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0196f
C14264 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# V_LOW 0.0113f
C14265 FULL_COUNTER.COUNT_SUB_DFF18.Q V_LOW 0.833f
C14266 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# sky130_fd_sc_hd__conb_1_40/HI 4.67e-19
C14267 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__conb_1_37/HI 0.00313f
C14268 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_1_107/Y 1.57e-20
C14269 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_7/LO 1.61e-21
C14270 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_47/a_791_47# 4.91e-20
C14271 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# V_GND 0.00385f
C14272 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__conb_1_29/LO 0.0134f
C14273 sky130_fd_sc_hd__inv_1_67/Y V_GND 1.37f
C14274 sky130_fd_sc_hd__conb_1_38/LO sky130_fd_sc_hd__inv_1_75/A 2.66e-21
C14275 sky130_fd_sc_hd__conb_1_13/LO V_GND -6.09e-19
C14276 sky130_fd_sc_hd__fill_8_819/VPB V_GND 0.408f
C14277 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 6.23e-19
C14278 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 3.01e-20
C14279 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.00133f
C14280 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# -4e-19
C14281 sky130_fd_sc_hd__dfbbn_1_29/a_1159_47# V_GND 0.00102f
C14282 sky130_fd_sc_hd__conb_1_30/LO RISING_COUNTER.COUNT_SUB_DFF5.Q 4.24e-19
C14283 sky130_fd_sc_hd__dfbbn_1_11/a_1340_413# V_GND 1.22e-19
C14284 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# V_LOW 0.0103f
C14285 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_68/A 0.00485f
C14286 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__conb_1_44/HI 0.01f
C14287 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.11e-19
C14288 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# V_LOW 0.00899f
C14289 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00168f
C14290 sky130_fd_sc_hd__dfbbn_1_8/a_581_47# V_GND -9.06e-19
C14291 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_36/LO 0.00525f
C14292 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# V_LOW -0.0119f
C14293 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 9.44e-20
C14294 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0674f
C14295 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 9.14e-19
C14296 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 9.68e-20
C14297 sky130_fd_sc_hd__dfbbn_1_36/a_1340_413# V_LOW -6.55e-19
C14298 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 2.93e-20
C14299 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# V_GND 0.00201f
C14300 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.69e-19
C14301 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0586f
C14302 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 1.28e-19
C14303 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0578f
C14304 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF0.Q 0.172f
C14305 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_45/LO 0.00572f
C14306 sky130_fd_sc_hd__inv_1_107/Y sky130_fd_sc_hd__conb_1_46/HI 0.0854f
C14307 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.22e-19
C14308 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# -2.57e-20
C14309 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 1.76e-19
C14310 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__inv_1_76/A 0.00142f
C14311 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_647_21# -0.00431f
C14312 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_473_413# -0.00461f
C14313 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 3.22e-21
C14314 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# Reset 0.00189f
C14315 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__inv_1_106/Y 1.19e-20
C14316 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 4.71e-20
C14317 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_791_47# 2.01e-20
C14318 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# V_GND 0.00165f
C14319 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 0.0427f
C14320 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# sky130_fd_sc_hd__conb_1_22/HI 2.07e-19
C14321 sky130_fd_sc_hd__inv_1_57/Y sky130_fd_sc_hd__conb_1_26/HI 0.309f
C14322 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# sky130_fd_sc_hd__inv_1_21/Y 9.65e-22
C14323 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# V_GND 5.9e-19
C14324 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF9.Q 8.97e-19
C14325 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# -0.00827f
C14326 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# -0.00117f
C14327 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# V_GND 1.65e-19
C14328 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0194f
C14329 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# V_LOW -0.107f
C14330 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 5.58e-19
C14331 sky130_fd_sc_hd__dfbbn_1_36/a_1159_47# V_GND -0.00168f
C14332 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_25/LO 9e-21
C14333 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# -0.00141f
C14334 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_43/HI 0.176f
C14335 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF11.Q 9.57e-20
C14336 Reset sky130_fd_sc_hd__inv_1_70/A 4.23e-20
C14337 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_19/Y 5.07e-22
C14338 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0497f
C14339 sky130_fd_sc_hd__conb_1_9/HI FULL_COUNTER.COUNT_SUB_DFF7.Q 0.13f
C14340 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0119f
C14341 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# sky130_fd_sc_hd__conb_1_27/HI 0.00447f
C14342 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# V_LOW -0.00722f
C14343 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# sky130_fd_sc_hd__inv_1_21/Y 0.00221f
C14344 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# -0.00813f
C14345 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0.00212f
C14346 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 0.00212f
C14347 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF4.Q 3.38e-21
C14348 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__conb_1_44/HI 0.0343f
C14349 sky130_fd_sc_hd__dfbbn_1_1/a_1340_413# V_LOW -6.55e-19
C14350 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# sky130_fd_sc_hd__conb_1_47/HI 0.00428f
C14351 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 0.0115f
C14352 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# V_LOW 0.00634f
C14353 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# sky130_fd_sc_hd__conb_1_47/HI -7.58e-20
C14354 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 0.017f
C14355 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# V_GND -0.00535f
C14356 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00143f
C14357 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__inv_1_12/Y 7.13e-22
C14358 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# sky130_fd_sc_hd__inv_1_65/Y 3.31e-19
C14359 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 3.87e-21
C14360 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 4.51e-19
C14361 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 6.87e-19
C14362 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__conb_1_13/HI 2.28e-19
C14363 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# sky130_fd_sc_hd__inv_1_12/Y 9.6e-20
C14364 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# V_GND 0.00208f
C14365 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__conb_1_24/HI 6.96e-20
C14366 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# -0.00141f
C14367 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 0.0142f
C14368 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_581_47# -2.6e-20
C14369 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 2.34e-19
C14370 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__inv_1_9/Y 7.13e-22
C14371 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 0.0569f
C14372 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# V_LOW 0.0122f
C14373 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00719f
C14374 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__conb_1_21/HI 5.47e-19
C14375 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0343f
C14376 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# V_LOW 1.79e-20
C14377 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.28f
C14378 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# sky130_fd_sc_hd__conb_1_37/HI 0.00836f
C14379 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# -3.79e-20
C14380 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1112_329# -0.00336f
C14381 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__inv_1_107/Y 2.27e-20
C14382 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 1.07e-19
C14383 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# sky130_fd_sc_hd__conb_1_32/HI 0.0169f
C14384 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00318f
C14385 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_20/Y 5.1e-19
C14386 sky130_fd_sc_hd__dfbbn_1_1/a_1159_47# V_GND 4.39e-19
C14387 sky130_fd_sc_hd__conb_1_18/LO FULL_COUNTER.COUNT_SUB_DFF5.Q 3.5e-21
C14388 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# V_LOW -0.0123f
C14389 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# sky130_fd_sc_hd__conb_1_29/LO 5.62e-20
C14390 sky130_fd_sc_hd__dfbbn_1_9/a_891_329# V_GND 4.61e-19
C14391 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__inv_16_1/Y 0.00384f
C14392 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__inv_1_71/A 4.43e-21
C14393 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__conb_1_34/HI 4.21e-20
C14394 sky130_fd_sc_hd__inv_1_50/Y V_GND 0.0432f
C14395 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 2.57e-19
C14396 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 6.05e-19
C14397 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 9.37e-21
C14398 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 3.25e-20
C14399 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# -2.32e-19
C14400 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -2.02e-19
C14401 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__conb_1_15/LO 0.00206f
C14402 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# V_LOW 1.79e-20
C14403 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__conb_1_36/LO 1.22e-20
C14404 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.19e-20
C14405 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# 0.00278f
C14406 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# V_LOW -0.00181f
C14407 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00256f
C14408 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# V_LOW -0.00663f
C14409 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_76/A 0.0532f
C14410 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.47e-20
C14411 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# V_GND -0.00709f
C14412 sky130_fd_sc_hd__inv_1_101/Y sky130_fd_sc_hd__conb_1_35/HI 3.47e-19
C14413 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__conb_1_13/HI 4.3e-19
C14414 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 3.59e-19
C14415 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# V_GND 1.64e-19
C14416 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 4.9e-21
C14417 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 5.72e-20
C14418 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_91/A 0.45f
C14419 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 3.24e-20
C14420 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 5.12e-20
C14421 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# V_GND -0.00515f
C14422 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# sky130_fd_sc_hd__conb_1_41/HI 1.06e-21
C14423 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.0029f
C14424 FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_16_1/Y 0.571f
C14425 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_193_47# -0.0146f
C14426 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00109f
C14427 sky130_fd_sc_hd__conb_1_50/LO V_GND -0.00279f
C14428 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.97e-21
C14429 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0153f
C14430 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# 0.0025f
C14431 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00182f
C14432 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_1_98/Y 5.73e-19
C14433 RISING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_28/HI 1.62e-19
C14434 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 2.84e-32
C14435 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_941_21# -1.62e-20
C14436 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# -2.32e-19
C14437 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0352f
C14438 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 0.0356f
C14439 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# V_LOW -9.94e-19
C14440 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# -4.5e-20
C14441 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# -1.64e-20
C14442 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.75e-20
C14443 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 9.87e-21
C14444 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 0.00105f
C14445 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 0.00142f
C14446 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 0.00599f
C14447 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0.00132f
C14448 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00237f
C14449 sky130_fd_sc_hd__dfbbn_1_10/Q_N FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00216f
C14450 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0.564f
C14451 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# -0.00117f
C14452 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# -0.00175f
C14453 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/a_941_21# -9.88e-20
C14454 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.3e-19
C14455 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.00163f
C14456 sky130_fd_sc_hd__dfbbn_1_41/Q_N sky130_fd_sc_hd__conb_1_27/HI -2.17e-19
C14457 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 1.13e-19
C14458 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# -0.00141f
C14459 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# sky130_fd_sc_hd__inv_1_21/Y 0.00371f
C14460 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_381_47# -0.00869f
C14461 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00278f
C14462 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_16/HI 3.05e-20
C14463 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_557_413# 3.12e-19
C14464 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 3.49e-20
C14465 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 3.49e-20
C14466 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 4.19e-20
C14467 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 7.63e-19
C14468 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 2.37e-19
C14469 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0965f
C14470 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 7.63e-19
C14471 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 2.37e-19
C14472 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0.00149f
C14473 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 1.71e-19
C14474 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 9.77e-19
C14475 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 1.01e-19
C14476 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__nand3_1_2/B 0.11f
C14477 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_43/a_791_47# 6.07e-20
C14478 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__inv_1_102/Y 3.94e-19
C14479 sky130_fd_sc_hd__dfbbn_1_40/Q_N sky130_fd_sc_hd__conb_1_47/HI -2.17e-19
C14480 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# sky130_fd_sc_hd__conb_1_36/HI 0.00217f
C14481 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# 0.0013f
C14482 sky130_fd_sc_hd__dfbbn_1_4/a_1363_47# V_GND 1.72e-19
C14483 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.79e-21
C14484 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 8.79e-22
C14485 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_48/Q_N 5.35e-19
C14486 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.0291f
C14487 sky130_fd_sc_hd__dfbbn_1_29/a_581_47# sky130_fd_sc_hd__inv_1_65/Y 5.8e-19
C14488 sky130_fd_sc_hd__nand2_8_3/Y sky130_fd_sc_hd__inv_1_67/Y 5.54e-19
C14489 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 0.0619f
C14490 sky130_fd_sc_hd__dfbbn_1_20/Q_N V_GND -0.00306f
C14491 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.77e-20
C14492 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 1.48e-20
C14493 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# V_LOW -0.00389f
C14494 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1159_47# 4e-20
C14495 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__conb_1_39/HI 1.05e-20
C14496 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 7.03e-20
C14497 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__conb_1_21/HI 3.23e-21
C14498 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# V_GND 3.4e-19
C14499 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/Q_N -4.78e-20
C14500 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_1_13/Y 1.63e-19
C14501 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_97/A 0.0156f
C14502 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_12/a_193_47# -4.7e-37
C14503 sky130_fd_sc_hd__dfbbn_1_23/a_1159_47# sky130_fd_sc_hd__conb_1_32/HI 0.00125f
C14504 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_16_2/Y 0.576f
C14505 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0162f
C14506 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0232f
C14507 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# V_LOW 1.79e-20
C14508 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__inv_1_15/Y 0.00498f
C14509 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__conb_1_2/LO 0.00638f
C14510 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_51/a_941_21# 3.56e-22
C14511 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# V_GND 0.0273f
C14512 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__conb_1_19/LO 1.33e-19
C14513 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__inv_1_15/Y 0.0401f
C14514 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0.00186f
C14515 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# -1.64e-19
C14516 FALLING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_103/Y 0.0277f
C14517 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 2.54e-20
C14518 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.39e-19
C14519 sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# V_GND 0.00116f
C14520 sky130_fd_sc_hd__conb_1_31/HI V_LOW 0.03f
C14521 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__conb_1_27/HI 2.53e-21
C14522 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# -3.72e-19
C14523 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# -0.00567f
C14524 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# V_LOW 0.0231f
C14525 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# V_GND -0.00815f
C14526 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.27e-19
C14527 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 2.31e-19
C14528 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0518f
C14529 sky130_fd_sc_hd__inv_1_56/Y sky130_fd_sc_hd__conb_1_26/HI 1.52e-20
C14530 sky130_fd_sc_hd__dfbbn_1_26/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00808f
C14531 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0101f
C14532 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0453f
C14533 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00598f
C14534 sky130_fd_sc_hd__inv_1_54/Y RISING_COUNTER.COUNT_SUB_DFF2.Q 0.407f
C14535 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 3e-21
C14536 sky130_fd_sc_hd__dfbbn_1_7/a_1363_47# V_GND -2.81e-19
C14537 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.73e-20
C14538 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1e-19
C14539 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 7.39e-20
C14540 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_17/HI 0.0577f
C14541 sky130_fd_sc_hd__inv_1_109/Y V_GND 0.0994f
C14542 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.138f
C14543 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00625f
C14544 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 0.00942f
C14545 sky130_fd_sc_hd__dfbbn_1_24/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.81e-19
C14546 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/Q_N 0.00975f
C14547 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 3.84e-20
C14548 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.00381f
C14549 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 0.0059f
C14550 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/Q_N -9.56e-20
C14551 sky130_fd_sc_hd__dfbbn_1_49/a_557_413# V_GND 3.03e-19
C14552 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# sky130_fd_sc_hd__conb_1_51/HI 0.00233f
C14553 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# sky130_fd_sc_hd__inv_1_76/A 0.00145f
C14554 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__inv_1_106/Y 0.00102f
C14555 sky130_fd_sc_hd__inv_1_68/A sky130_fd_sc_hd__inv_1_70/A 0.387f
C14556 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 1.4e-20
C14557 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 2.39e-20
C14558 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0.00893f
C14559 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 2.41e-19
C14560 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# V_LOW 0.0303f
C14561 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.79e-21
C14562 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_89/Y 4.56e-21
C14563 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__conb_1_33/LO 0.0537f
C14564 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 5.2e-19
C14565 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 4.46e-21
C14566 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__conb_1_23/HI 4.7e-20
C14567 sky130_fd_sc_hd__dfbbn_1_38/Q_N FALLING_COUNTER.COUNT_SUB_DFF10.Q 2.34e-19
C14568 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 6.69e-20
C14569 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0.00128f
C14570 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.16e-21
C14571 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00399f
C14572 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# -0.00107f
C14573 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.45e-19
C14574 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# V_LOW -0.00121f
C14575 sky130_fd_sc_hd__conb_1_27/HI Reset 1.41e-19
C14576 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 2.27e-20
C14577 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00174f
C14578 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 2.27e-20
C14579 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_43/A 0.0255f
C14580 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_557_413# -3.67e-20
C14581 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# -0.00381f
C14582 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_21/HI 6.28e-20
C14583 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__inv_1_102/Y 8.82e-20
C14584 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__conb_1_4/LO 0.0116f
C14585 sky130_fd_sc_hd__conb_1_45/HI V_GND 0.198f
C14586 sky130_fd_sc_hd__dfbbn_1_9/Q_N V_LOW -0.00253f
C14587 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# V_LOW -4.1e-19
C14588 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# sky130_fd_sc_hd__conb_1_36/HI 6.97e-20
C14589 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__inv_1_8/Y 0.0107f
C14590 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# V_LOW 3.56e-20
C14591 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_41/LO 0.00904f
C14592 sky130_fd_sc_hd__inv_1_53/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 2.73e-20
C14593 sky130_fd_sc_hd__dfbbn_1_17/a_557_413# V_GND 2.63e-19
C14594 sky130_fd_sc_hd__nand2_8_4/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00464f
C14595 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# 2.52e-19
C14596 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.1e-19
C14597 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 1.07e-20
C14598 FALLING_COUNTER.COUNT_SUB_DFF11.Q V_GND 3.23f
C14599 sky130_fd_sc_hd__inv_1_43/A sky130_fd_sc_hd__inv_1_45/A 0.00226f
C14600 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.17e-19
C14601 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# sky130_fd_sc_hd__conb_1_41/HI -2.65e-20
C14602 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__inv_1_90/Y 4.23e-21
C14603 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 1.04e-19
C14604 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 2.86e-20
C14605 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 9.57e-21
C14606 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# V_GND -0.00463f
C14607 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 5.98e-19
C14608 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 3.34e-19
C14609 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 2.75e-19
C14610 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0.00159f
C14611 sky130_fd_sc_hd__inv_1_89/A sky130_fd_sc_hd__inv_1_83/Y 0.0362f
C14612 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0312f
C14613 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.144f
C14614 FALLING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__inv_1_106/Y 0.00334f
C14615 sky130_fd_sc_hd__dfbbn_1_43/a_891_329# V_GND 3.7e-19
C14616 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_193_47# -0.179f
C14617 sky130_fd_sc_hd__conb_1_20/HI CLOCK_GEN.SR_Op.Q 1.15e-19
C14618 sky130_fd_sc_hd__dfbbn_1_3/a_1340_413# V_GND 1.64e-19
C14619 sky130_fd_sc_hd__conb_1_21/LO sky130_fd_sc_hd__conb_1_21/HI 0.00889f
C14620 sky130_fd_sc_hd__dfbbn_1_39/Q_N FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.24e-19
C14621 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__inv_16_1/Y 0.0618f
C14622 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# sky130_fd_sc_hd__inv_1_15/Y 0.00104f
C14623 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__inv_1_16/Y 7.25e-19
C14624 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 1.65e-19
C14625 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00102f
C14626 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__conb_1_12/HI 6.6e-19
C14627 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# -1.66e-19
C14628 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# V_LOW 0.00983f
C14629 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 6.77e-20
C14630 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__conb_1_16/LO 1.38e-19
C14631 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# -2.37e-19
C14632 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -0.013f
C14633 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 3.53e-19
C14634 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_47/Y 0.0708f
C14635 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# sky130_fd_sc_hd__conb_1_32/HI 2.12e-21
C14636 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0.00502f
C14637 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0308f
C14638 sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__inv_1_27/Y 0.0409f
C14639 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_32/Y 5.47e-20
C14640 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_34/A 0.011f
C14641 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__conb_1_35/HI 0.014f
C14642 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 1.02e-19
C14643 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 0.0265f
C14644 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 1.95e-20
C14645 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0138f
C14646 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.0132f
C14647 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# 0.00255f
C14648 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# 2.06e-20
C14649 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 0.00429f
C14650 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 4.06e-21
C14651 RISING_COUNTER.COUNT_SUB_DFF6.Q V_GND 4.58f
C14652 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00515f
C14653 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.71e-20
C14654 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__conb_1_46/HI 0.00386f
C14655 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0275f
C14656 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/Q_N -9.56e-20
C14657 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.12e-19
C14658 sky130_fd_sc_hd__conb_1_10/LO sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 7.06e-20
C14659 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 8.12e-19
C14660 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 9.78e-19
C14661 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 7.19e-19
C14662 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# V_LOW 0.0066f
C14663 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_16_2/Y 0.216f
C14664 sky130_fd_sc_hd__inv_1_97/A sky130_fd_sc_hd__inv_1_86/Y 0.0915f
C14665 sky130_fd_sc_hd__inv_1_39/A V_GND 0.105f
C14666 sky130_fd_sc_hd__inv_1_76/A sky130_fd_sc_hd__inv_2_0/Y 0.0425f
C14667 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00509f
C14668 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_16_1/Y 0.00142f
C14669 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 0.00881f
C14670 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_791_47# 3.3e-21
C14671 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 0.00387f
C14672 sky130_fd_sc_hd__conb_1_27/HI sky130_fd_sc_hd__inv_1_57/Y 2.04e-20
C14673 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00631f
C14674 sky130_fd_sc_hd__dfbbn_1_8/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 2.91e-19
C14675 sky130_fd_sc_hd__conb_1_43/LO sky130_fd_sc_hd__inv_1_105/Y 0.0107f
C14676 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 6.4e-19
C14677 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__conb_1_33/HI 0.0124f
C14678 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__conb_1_46/HI 0.0181f
C14679 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__nand2_8_2/A 0.0558f
C14680 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# sky130_fd_sc_hd__conb_1_2/HI 8.64e-19
C14681 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.0139f
C14682 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# -0.0586f
C14683 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# -4.36e-19
C14684 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 5.52e-20
C14685 sky130_fd_sc_hd__conb_1_15/HI V_LOW 0.188f
C14686 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# sky130_fd_sc_hd__conb_1_47/HI 5.06e-20
C14687 sky130_fd_sc_hd__inv_1_90/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 4.56e-21
C14688 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 2.02e-19
C14689 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0272f
C14690 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.78e-19
C14691 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 6.61e-20
C14692 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 5.64e-20
C14693 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 5.52e-19
C14694 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# 8.91e-21
C14695 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 6.1e-19
C14696 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__conb_1_45/HI 0.0157f
C14697 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# V_LOW 0.0161f
C14698 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# V_LOW 0.00769f
C14699 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 0.0019f
C14700 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0235f
C14701 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 7.16e-20
C14702 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 1.47e-21
C14703 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_21/HI 0.0259f
C14704 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# V_LOW 0.0053f
C14705 sky130_fd_sc_hd__conb_1_14/LO sky130_fd_sc_hd__inv_16_2/Y 4.88e-20
C14706 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# V_LOW 0.028f
C14707 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 7.24e-19
C14708 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0366f
C14709 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_1_13/Y 7.33e-20
C14710 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 0.0301f
C14711 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# V_LOW 9.19e-19
C14712 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0373f
C14713 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.97e-20
C14714 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 0.00198f
C14715 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.00344f
C14716 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 0.0122f
C14717 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 4.76e-19
C14718 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 4.03e-19
C14719 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 4.03e-19
C14720 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 4.76e-19
C14721 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 0.00865f
C14722 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# V_LOW 0.0139f
C14723 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_119/Y 0.0169f
C14724 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# V_GND -2.59e-19
C14725 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# V_GND -0.00364f
C14726 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__conb_1_22/HI 3.13e-19
C14727 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 0.0298f
C14728 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_647_21# -6.43e-20
C14729 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_473_413# -3.06e-20
C14730 sky130_fd_sc_hd__dfbbn_1_15/a_891_329# V_GND 4.09e-19
C14731 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.00477f
C14732 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# V_GND 0.00393f
C14733 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# -7.17e-20
C14734 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# -1.66e-19
C14735 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 1.22e-20
C14736 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# 0.00136f
C14737 FALLING_COUNTER.COUNT_SUB_DFF5.Q V_LOW 1.9f
C14738 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 0.00145f
C14739 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# V_GND -0.00658f
C14740 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__conb_1_35/HI 2.59e-19
C14741 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__inv_1_76/A 1.74e-19
C14742 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/Q_N 4.53e-21
C14743 sky130_fd_sc_hd__nor2_1_0/a_109_297# V_GND -9.61e-19
C14744 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# sky130_fd_sc_hd__inv_16_1/Y 1.15e-19
C14745 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# 1.29e-20
C14746 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 1.33e-19
C14747 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 8.49e-20
C14748 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.52e-19
C14749 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_40/HI 4.15e-20
C14750 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 0.124f
C14751 sky130_fd_sc_hd__dfbbn_1_51/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0139f
C14752 RISING_COUNTER.COUNT_SUB_DFF1.Q RISING_COUNTER.COUNT_SUB_DFF2.Q 2.53f
C14753 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_11/HI 7.49e-20
C14754 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF9.Q 3.02e-19
C14755 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__conb_1_49/HI 5.09e-19
C14756 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__inv_1_106/Y 0.0123f
C14757 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# V_GND -0.00398f
C14758 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__inv_1_15/Y 0.0163f
C14759 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_45/LO 0.0453f
C14760 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_59/Y 0.21f
C14761 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_63/Y 4.38e-20
C14762 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# V_GND 0.00436f
C14763 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0402f
C14764 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0386f
C14765 sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.3e-20
C14766 sky130_fd_sc_hd__inv_1_19/Y V_LOW 0.198f
C14767 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_11/Y 0.0557f
C14768 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00172f
C14769 FULL_COUNTER.COUNT_SUB_DFF19.Q CLOCK_GEN.SR_Op.Q 5.2e-20
C14770 sky130_fd_sc_hd__dfbbn_1_17/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.48e-19
C14771 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 0.0136f
C14772 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# V_LOW 0.00715f
C14773 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 0.0012f
C14774 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0381f
C14775 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_0/HI 0.293f
C14776 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# sky130_fd_sc_hd__inv_1_23/Y 0.0191f
C14777 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 0.00132f
C14778 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 6.97e-22
C14779 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_43/HI 0.0832f
C14780 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# sky130_fd_sc_hd__conb_1_46/HI 0.0069f
C14781 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_95/A 0.00492f
C14782 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.91e-19
C14783 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_50/A 0.00114f
C14784 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_43/A 0.00326f
C14785 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# sky130_fd_sc_hd__inv_1_21/Y 4.67e-19
C14786 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 6.64e-21
C14787 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__inv_16_2/Y 0.0495f
C14788 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__inv_1_20/Y 0.0107f
C14789 sky130_fd_sc_hd__dfbbn_1_43/Q_N V_LOW -0.00141f
C14790 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF9.Q 3e-21
C14791 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_62/Y 0.124f
C14792 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# -5.72e-19
C14793 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# -0.0103f
C14794 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# V_GND -0.00169f
C14795 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__inv_1_11/Y 4.98e-19
C14796 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF18.Q 4.75e-20
C14797 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.79e-19
C14798 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 3.53e-20
C14799 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 1.27e-20
C14800 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.34e-19
C14801 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.67e-19
C14802 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_37/a_1363_47# 3.91e-19
C14803 sky130_fd_sc_hd__dfbbn_1_26/a_1340_413# V_LOW -6.55e-19
C14804 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.4e-19
C14805 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 3.4e-20
C14806 sky130_fd_sc_hd__conb_1_21/LO CLOCK_GEN.SR_Op.Q 0.0324f
C14807 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_1_17/Y 0.0188f
C14808 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# V_LOW 1.73e-20
C14809 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 9.59e-19
C14810 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 4.82e-21
C14811 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.58e-20
C14812 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# V_LOW 2.94e-20
C14813 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_67/Y 5.59e-21
C14814 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__dfbbn_1_13/a_1112_329# -0.00336f
C14815 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/Q_N 1.39e-19
C14816 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# sky130_fd_sc_hd__inv_1_100/Y 0.00813f
C14817 sky130_fd_sc_hd__dfbbn_1_13/a_581_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.79e-19
C14818 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.016f
C14819 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# V_LOW -2.94e-19
C14820 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.35e-21
C14821 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__conb_1_46/HI 3.49e-21
C14822 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 5.54e-20
C14823 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__conb_1_50/LO 6.57e-20
C14824 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00104f
C14825 sky130_fd_sc_hd__inv_1_89/A V_LOW 0.195f
C14826 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 7.64e-19
C14827 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0.00131f
C14828 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 0.00131f
C14829 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 7.64e-19
C14830 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__inv_1_17/Y 2.97e-19
C14831 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 6.14e-21
C14832 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# V_GND 0.00625f
C14833 sky130_fd_sc_hd__dfbbn_1_26/a_1159_47# V_GND -0.00156f
C14834 sky130_fd_sc_hd__dfbbn_1_44/a_1112_329# V_LOW 4.8e-20
C14835 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# sky130_fd_sc_hd__inv_1_105/Y 0.00215f
C14836 sky130_fd_sc_hd__dfbbn_1_4/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 0.00105f
C14837 sky130_fd_sc_hd__dfbbn_1_31/a_1159_47# V_GND 6.11e-19
C14838 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_1_75/Y 5.46e-20
C14839 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.36e-19
C14840 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# 4.06e-21
C14841 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# V_GND -0.0152f
C14842 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__dfbbn_1_14/Q_N 0.00133f
C14843 sky130_fd_sc_hd__conb_1_46/LO FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0104f
C14844 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__conb_1_35/HI 6.62e-19
C14845 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# V_LOW 0.00665f
C14846 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# CLOCK_GEN.SR_Op.Q 2.09e-19
C14847 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 8.21e-19
C14848 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# V_GND 0.00388f
C14849 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_891_329# -2.2e-20
C14850 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# -0.00106f
C14851 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__conb_1_46/HI 1.55e-20
C14852 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0113f
C14853 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_891_329# -2.2e-20
C14854 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# -0.00161f
C14855 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.01e-20
C14856 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.29e-20
C14857 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 3.5e-22
C14858 sky130_fd_sc_hd__inv_1_96/A sky130_fd_sc_hd__inv_1_71/Y 2.88e-20
C14859 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__inv_1_106/Y 0.0117f
C14860 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# V_GND -0.0128f
C14861 sky130_fd_sc_hd__dfbbn_1_44/a_581_47# V_GND 2.66e-19
C14862 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 4.56e-21
C14863 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.00427f
C14864 FALLING_COUNTER.COUNT_SUB_DFF8.Q V_GND 0.594f
C14865 sky130_fd_sc_hd__conb_1_2/HI sky130_fd_sc_hd__inv_16_2/Y 0.0909f
C14866 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0536f
C14867 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__conb_1_42/HI 4.88e-19
C14868 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 4.07e-20
C14869 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_1_5/Y 1.53e-19
C14870 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00364f
C14871 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 1.62e-19
C14872 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.17e-22
C14873 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 5.16e-20
C14874 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0295f
C14875 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -0.00395f
C14876 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# -0.0158f
C14877 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 5.4e-19
C14878 sky130_fd_sc_hd__dfbbn_1_51/a_891_329# V_GND 3.46e-19
C14879 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 1.09e-19
C14880 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# sky130_fd_sc_hd__inv_1_23/Y 0.0505f
C14881 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# -9.88e-20
C14882 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# -6.23e-21
C14883 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# -0.00175f
C14884 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0177f
C14885 FALLING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_106/Y 0.0339f
C14886 sky130_fd_sc_hd__inv_1_99/Y sky130_fd_sc_hd__inv_1_108/Y 3.03e-19
C14887 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 2.1e-20
C14888 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.14e-21
C14889 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__inv_1_10/Y 0.00132f
C14890 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.93e-21
C14891 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__nand2_8_9/Y 3.68e-21
C14892 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.00166f
C14893 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 0.00166f
C14894 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00775f
C14895 sky130_fd_sc_hd__dfbbn_1_39/Q_N sky130_fd_sc_hd__conb_1_46/HI -2.17e-19
C14896 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0.00946f
C14897 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_42/a_381_47# -3.79e-20
C14898 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_42/a_1112_329# -4.66e-20
C14899 sky130_fd_sc_hd__dfbbn_1_7/a_1159_47# sky130_fd_sc_hd__inv_16_2/Y 0.00138f
C14900 FALLING_COUNTER.COUNT_SUB_DFF15.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0206f
C14901 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# sky130_fd_sc_hd__conb_1_2/HI 4.96e-19
C14902 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 1.32e-20
C14903 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_16_0/Y 0.507f
C14904 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_63/Y 5.95e-19
C14905 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# -1.24e-20
C14906 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__inv_1_54/Y 7.96e-19
C14907 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__inv_1_11/Y 1.21e-19
C14908 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__dfbbn_1_23/a_1340_413# -6.8e-19
C14909 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00215f
C14910 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_1_60/Y 6.78e-19
C14911 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# V_GND -0.00177f
C14912 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# sky130_fd_sc_hd__inv_1_11/Y 8.03e-21
C14913 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__inv_1_54/Y 1.4e-21
C14914 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -0.00746f
C14915 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_473_413# -0.00563f
C14916 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.34e-19
C14917 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.366f
C14918 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0037f
C14919 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__conb_1_9/HI 6.82e-20
C14920 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/Q_N 7.72e-21
C14921 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# -6.43e-19
C14922 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_473_413# -0.0225f
C14923 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.067f
C14924 sky130_fd_sc_hd__dfbbn_1_15/Q_N V_LOW 0.00119f
C14925 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# V_LOW -0.113f
C14926 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 4.43e-21
C14927 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 2.7e-21
C14928 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 5.14e-20
C14929 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 9.88e-19
C14930 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 9.77e-19
C14931 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 1.84e-20
C14932 sky130_fd_sc_hd__conb_1_48/HI V_LOW 0.0124f
C14933 sky130_fd_sc_hd__nand2_8_0/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 0.00329f
C14934 sky130_fd_sc_hd__dfbbn_1_19/a_1340_413# V_LOW -6.55e-19
C14935 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__inv_1_5/Y 8.81e-19
C14936 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 2.34e-20
C14937 sky130_fd_sc_hd__dfbbn_1_31/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.00202f
C14938 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# sky130_fd_sc_hd__conb_1_25/HI 0.0137f
C14939 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__inv_1_90/Y 0.0704f
C14940 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# sky130_fd_sc_hd__inv_1_17/Y 4.98e-21
C14941 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 3.52e-19
C14942 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.1e-20
C14943 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# V_GND -0.00509f
C14944 sky130_fd_sc_hd__dfbbn_1_27/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 8.13e-21
C14945 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.346f
C14946 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -6.23e-21
C14947 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# -0.00527f
C14948 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# V_LOW -0.107f
C14949 FULL_COUNTER.COUNT_SUB_DFF16.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0263f
C14950 sky130_fd_sc_hd__conb_1_38/HI FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.465f
C14951 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.00219f
C14952 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_581_47# 1.02e-19
C14953 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 2.48e-20
C14954 sky130_fd_sc_hd__dfbbn_1_19/a_1159_47# V_GND 3.92e-19
C14955 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# -0.00376f
C14956 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# sky130_fd_sc_hd__inv_16_0/Y 0.0012f
C14957 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_25/a_381_47# 1.34e-19
C14958 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__inv_1_47/Y 2.41e-19
C14959 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# sky130_fd_sc_hd__inv_16_1/Y 1.31e-19
C14960 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 1.51e-21
C14961 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 5.99e-19
C14962 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 2.83e-19
C14963 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0163f
C14964 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# -3.46e-20
C14965 sky130_fd_sc_hd__inv_1_98/Y sky130_fd_sc_hd__conb_1_37/HI 0.0271f
C14966 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 2.62e-20
C14967 sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 4.04e-20
C14968 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_381_47# -0.00813f
C14969 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 1.53e-19
C14970 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# sky130_fd_sc_hd__inv_1_19/Y 0.022f
C14971 sky130_fd_sc_hd__conb_1_41/LO FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.00659f
C14972 sky130_fd_sc_hd__conb_1_38/HI V_LOW 0.195f
C14973 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 0.00518f
C14974 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 0.0289f
C14975 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF4.Q 1.6e-19
C14976 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# Reset 1.6e-19
C14977 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 3.23e-21
C14978 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 6.31e-21
C14979 sky130_fd_sc_hd__inv_1_1/Y V_GND 0.0433f
C14980 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__conb_1_23/HI 1.52e-20
C14981 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__inv_1_11/Y 6.42e-20
C14982 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# V_GND 0.00402f
C14983 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# sky130_fd_sc_hd__conb_1_29/LO 8.84e-20
C14984 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_1340_413# -6.8e-19
C14985 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 2.3e-22
C14986 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0108f
C14987 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__conb_1_20/HI 2.75e-19
C14988 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 5.13e-21
C14989 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_112/Y 0.00446f
C14990 sky130_fd_sc_hd__dfbbn_1_5/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF11.Q 1.71e-21
C14991 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 3.58e-19
C14992 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 1.57e-20
C14993 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 6.08e-20
C14994 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 4.29e-19
C14995 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 6.08e-20
C14996 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 4.29e-19
C14997 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__inv_16_2/Y 0.104f
C14998 sky130_fd_sc_hd__inv_1_7/Y FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0122f
C14999 sky130_fd_sc_hd__conb_1_23/LO RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0766f
C15000 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# -5.33e-20
C15001 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_557_413# -3.67e-20
C15002 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# CLOCK_GEN.SR_Op.Q 5.63e-19
C15003 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 1.41e-19
C15004 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__inv_1_20/Y 1.63e-20
C15005 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 7.53e-21
C15006 RISING_COUNTER.COUNT_SUB_DFF0.Q RISING_COUNTER.COUNT_SUB_DFF11.Q 2.75e-19
C15007 sky130_fd_sc_hd__conb_1_7/LO FULL_COUNTER.COUNT_SUB_DFF9.Q 3.25e-19
C15008 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0.00113f
C15009 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00132f
C15010 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_581_47# -2.6e-20
C15011 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# sky130_fd_sc_hd__inv_1_60/Y 4.61e-19
C15012 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 0.0107f
C15013 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# -9.41e-19
C15014 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# sky130_fd_sc_hd__inv_1_55/Y 1.32e-21
C15015 sky130_fd_sc_hd__dfbbn_1_30/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 2.66e-20
C15016 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# V_LOW 0.00207f
C15017 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0116f
C15018 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_381_47# 0.00146f
C15019 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# -6.8e-19
C15020 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0428f
C15021 sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# V_LOW -2.68e-19
C15022 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# sky130_fd_sc_hd__inv_16_0/Y 2.34e-19
C15023 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 0.00617f
C15024 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__conb_1_6/HI 0.025f
C15025 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 1.51e-19
C15026 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 1.06e-19
C15027 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 1.18e-21
C15028 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.16e-19
C15029 sky130_fd_sc_hd__dfbbn_1_0/a_581_47# sky130_fd_sc_hd__inv_1_5/Y 2.34e-19
C15030 sky130_fd_sc_hd__conb_1_12/HI V_LOW 0.155f
C15031 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 1.23e-20
C15032 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand3_1_2/Y 0.00445f
C15033 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 6.98e-20
C15034 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__conb_1_48/HI 0.0056f
C15035 sky130_fd_sc_hd__conb_1_12/HI sky130_fd_sc_hd__conb_1_13/HI 5.61e-21
C15036 sky130_fd_sc_hd__inv_1_97/A V_GND 0.241f
C15037 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# sky130_fd_sc_hd__inv_1_9/Y 2.63e-19
C15038 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# V_GND -5.53e-19
C15039 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.57e-19
C15040 sky130_fd_sc_hd__dfbbn_1_30/a_1363_47# V_GND 1.64e-19
C15041 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 2.57e-20
C15042 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0794f
C15043 sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 0.00151f
C15044 sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# V_LOW -2.68e-19
C15045 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0011f
C15046 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/Q_N -6.48e-19
C15047 FALLING_COUNTER.COUNT_SUB_DFF13.Q V_GND 0.699f
C15048 sky130_fd_sc_hd__dfbbn_1_51/Q_N V_LOW 6.79e-19
C15049 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_891_329# 1.48e-20
C15050 sky130_fd_sc_hd__nand2_1_5/Y V_LOW 0.0152f
C15051 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00806f
C15052 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_13/Y 3.07e-21
C15053 sky130_fd_sc_hd__dfbbn_1_40/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 8.14e-20
C15054 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 9.08e-21
C15055 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 1.2e-21
C15056 sky130_fd_sc_hd__dfbbn_1_2/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0188f
C15057 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# sky130_fd_sc_hd__conb_1_24/HI 7.11e-21
C15058 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# V_GND 0.062f
C15059 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 1.02e-19
C15060 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 9.59e-19
C15061 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# -0.00107f
C15062 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_1_48/Y 0.136f
C15063 FULL_COUNTER.COUNT_SUB_DFF6.Q FULL_COUNTER.COUNT_SUB_DFF7.Q 0.526f
C15064 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 8.73e-21
C15065 sky130_fd_sc_hd__conb_1_18/HI V_LOW 0.121f
C15066 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 1.67e-20
C15067 sky130_fd_sc_hd__inv_1_119/Y transmission_gate_0/GN 0.0254f
C15068 sky130_fd_sc_hd__nand2_8_1/a_27_47# sky130_fd_sc_hd__nand3_1_2/B 0.061f
C15069 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 0.00578f
C15070 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 5.82e-19
C15071 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0299f
C15072 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__conb_1_5/HI 2.27e-19
C15073 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_27/HI 0.0012f
C15074 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# V_GND 1.75e-19
C15075 sky130_fd_sc_hd__inv_1_18/Y V_GND 0.0902f
C15076 sky130_fd_sc_hd__conb_1_30/HI sky130_fd_sc_hd__conb_1_22/HI 2.52e-20
C15077 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 2.91e-21
C15078 sky130_fd_sc_hd__dfbbn_1_13/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0315f
C15079 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__conb_1_28/HI 0.00726f
C15080 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# sky130_fd_sc_hd__conb_1_20/HI -2.65e-20
C15081 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0446f
C15082 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# sky130_fd_sc_hd__inv_1_8/Y 7.42e-20
C15083 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_50/A 7.58e-19
C15084 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 3.04e-20
C15085 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 6.8e-20
C15086 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 5.47e-20
C15087 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__dfbbn_1_26/Q_N 5.47e-20
C15088 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_2/A 0.152f
C15089 sky130_fd_sc_hd__nand2_8_3/A V_GND 0.049f
C15090 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_26/LO 6.88e-19
C15091 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__conb_1_44/HI 6.96e-22
C15092 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF7.Q 1.27e-19
C15093 sky130_fd_sc_hd__dfbbn_1_3/Q_N sky130_fd_sc_hd__conb_1_2/HI 0.00667f
C15094 sky130_fd_sc_hd__fill_4_63/VPB V_LOW 0.797f
C15095 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 4.36e-19
C15096 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 4.3e-19
C15097 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 3.04e-19
C15098 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.65e-20
C15099 sky130_fd_sc_hd__conb_1_31/LO sky130_fd_sc_hd__inv_1_62/Y 0.0844f
C15100 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__inv_1_58/Y 1.77e-19
C15101 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__conb_1_23/HI -0.00192f
C15102 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# sky130_fd_sc_hd__inv_16_2/Y 0.00526f
C15103 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 1.89e-20
C15104 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.74e-19
C15105 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 2.99e-20
C15106 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 3.42e-19
C15107 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 3.55e-21
C15108 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# sky130_fd_sc_hd__conb_1_25/HI 0.00929f
C15109 FULL_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_15/Y 7.76e-20
C15110 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 3.37e-19
C15111 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0373f
C15112 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_31/HI 0.00291f
C15113 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.62e-19
C15114 sky130_fd_sc_hd__conb_1_13/LO sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 4.7e-21
C15115 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__conb_1_16/LO 0.0618f
C15116 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# sky130_fd_sc_hd__inv_1_101/Y 0.00157f
C15117 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0211f
C15118 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_40/HI 0.00188f
C15119 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 2.75e-20
C15120 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.00755f
C15121 sky130_fd_sc_hd__dfbbn_1_43/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.24e-19
C15122 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_97/Y 4.71e-19
C15123 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# CLOCK_GEN.SR_Op.Q 0.00212f
C15124 sky130_fd_sc_hd__dfbbn_1_21/a_557_413# V_LOW -9.15e-19
C15125 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF4.Q 2.55e-19
C15126 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# FULL_COUNTER.COUNT_SUB_DFF10.Q 5.67e-19
C15127 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# V_GND 0.00635f
C15128 sky130_fd_sc_hd__conb_1_0/HI FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00286f
C15129 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_1_105/Y 0.00133f
C15130 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_78/A 0.0512f
C15131 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# sky130_fd_sc_hd__inv_1_54/Y 0.00548f
C15132 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__conb_1_2/HI 0.0699f
C15133 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.71e-19
C15134 sky130_fd_sc_hd__conb_1_24/HI RISING_COUNTER.COUNT_SUB_DFF4.Q 4.91e-19
C15135 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 5.74e-19
C15136 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 5.82e-20
C15137 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 4.39e-19
C15138 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.0036f
C15139 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 9.65e-21
C15140 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.13e-21
C15141 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 0.422f
C15142 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# sky130_fd_sc_hd__inv_1_11/Y 7.8e-22
C15143 sky130_fd_sc_hd__dfbbn_1_41/Q_N RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0299f
C15144 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# sky130_fd_sc_hd__inv_16_0/Y 4.76e-19
C15145 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 8.31e-20
C15146 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 7.32e-20
C15147 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.14e-19
C15148 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_76/A 0.069f
C15149 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__inv_1_18/Y 1.56e-19
C15150 sky130_fd_sc_hd__conb_1_9/HI V_LOW 0.0333f
C15151 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_16_1/Y 0.00855f
C15152 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# sky130_fd_sc_hd__conb_1_6/HI 3.15e-21
C15153 sky130_fd_sc_hd__dfbbn_1_21/a_1340_413# V_GND 1.26e-19
C15154 sky130_fd_sc_hd__inv_1_61/Y RISING_COUNTER.COUNT_SUB_DFF4.Q 1.31e-20
C15155 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__inv_1_68/A 0.0203f
C15156 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0619f
C15157 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 0.574f
C15158 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__inv_1_112/Y 7.9e-21
C15159 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 4.57e-22
C15160 sky130_fd_sc_hd__conb_1_16/HI V_GND 0.148f
C15161 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# sky130_fd_sc_hd__conb_1_42/HI 7.74e-20
C15162 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__conb_1_22/HI 1.61e-20
C15163 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0201f
C15164 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_381_47# 1.9e-19
C15165 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# V_GND 0.0105f
C15166 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.61e-19
C15167 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0399f
C15168 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.0125f
C15169 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__inv_1_99/Y 0.00382f
C15170 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 2.32e-19
C15171 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__conb_1_28/HI 0.00971f
C15172 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0155f
C15173 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0.00283f
C15174 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0.00277f
C15175 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 2.15e-19
C15176 sky130_fd_sc_hd__conb_1_12/LO V_LOW 0.0672f
C15177 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 1.55e-20
C15178 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_50/a_193_47# 2.95e-19
C15179 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 4.04e-21
C15180 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_473_413# -0.0222f
C15181 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# -0.0114f
C15182 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_381_47# -2.53e-20
C15183 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_6/Y 0.0239f
C15184 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 1.12f
C15185 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__conb_1_44/HI 3.97e-20
C15186 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.62e-20
C15187 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0351f
C15188 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_18/HI 3.27e-19
C15189 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# sky130_fd_sc_hd__inv_1_98/Y 3.82e-19
C15190 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__nand2_1_5/a_113_47# 4.44e-20
C15191 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# V_GND 0.0127f
C15192 sky130_fd_sc_hd__inv_1_93/Y sky130_fd_sc_hd__inv_1_97/Y 8.18e-20
C15193 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# sky130_fd_sc_hd__conb_1_18/HI -1.88e-20
C15194 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__nand2_1_0/Y 7.76e-19
C15195 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_17/HI 4.91e-21
C15196 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__conb_1_32/HI 0.0446f
C15197 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00224f
C15198 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# sky130_fd_sc_hd__inv_16_2/Y 0.0402f
C15199 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.46e-19
C15200 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 5.74e-20
C15201 sky130_fd_sc_hd__dfbbn_1_20/Q_N sky130_fd_sc_hd__inv_1_55/Y 4.84e-20
C15202 sky130_fd_sc_hd__conb_1_9/LO V_GND -0.00315f
C15203 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 0.00471f
C15204 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# 4.88e-19
C15205 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.2e-20
C15206 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_193_47# -0.0175f
C15207 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 0.0108f
C15208 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF13.Q 3.5e-19
C15209 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# sky130_fd_sc_hd__conb_1_30/HI 4.94e-19
C15210 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# -0.00615f
C15211 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_557_413# -3.67e-20
C15212 sky130_fd_sc_hd__dfbbn_1_9/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 3.04e-19
C15213 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 5.46e-20
C15214 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_95/A 0.0124f
C15215 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_647_21# 0.0261f
C15216 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 8.83e-22
C15217 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 2.97e-20
C15218 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 1.18e-20
C15219 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 1.06e-21
C15220 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__conb_1_18/HI 1.82e-19
C15221 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# sky130_fd_sc_hd__conb_1_22/HI 0.0446f
C15222 sky130_fd_sc_hd__dfbbn_1_7/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF17.Q 5.37e-20
C15223 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_193_47# -0.154f
C15224 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 1.71e-19
C15225 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 5.29e-20
C15226 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_18/Y 2.26e-20
C15227 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__conb_1_39/HI 8.45e-19
C15228 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# sky130_fd_sc_hd__conb_1_16/HI 0.012f
C15229 RISING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_22/HI 0.536f
C15230 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__nand2_8_9/Y 5.67e-20
C15231 sky130_fd_sc_hd__dfbbn_1_37/a_557_413# V_LOW 3.56e-20
C15232 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00223f
C15233 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# V_LOW 0.0131f
C15234 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_647_21# 4.65e-19
C15235 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__conb_1_12/HI -0.00239f
C15236 sky130_fd_sc_hd__inv_1_62/Y V_LOW 0.106f
C15237 sky130_fd_sc_hd__dfbbn_1_48/a_581_47# sky130_fd_sc_hd__inv_16_0/Y 3.49e-20
C15238 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 1.45e-20
C15239 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 3.49e-21
C15240 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 1.72e-20
C15241 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__inv_1_102/Y 2.61e-20
C15242 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# V_LOW -0.113f
C15243 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_381_47# -0.00144f
C15244 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0014f
C15245 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0274f
C15246 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# sky130_fd_sc_hd__conb_1_6/HI 3.08e-21
C15247 Reset RISING_COUNTER.COUNT_SUB_DFF3.Q 3.03e-19
C15248 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_26/HI 7.14e-20
C15249 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_76/A 7.33e-19
C15250 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00104f
C15251 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.016f
C15252 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0193f
C15253 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1112_329# 0.00226f
C15254 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF14.Q 1e-19
C15255 sky130_fd_sc_hd__conb_1_21/HI V_GND 0.0659f
C15256 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__inv_1_23/Y 0.00667f
C15257 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# -0.0128f
C15258 sky130_fd_sc_hd__conb_1_8/HI FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0418f
C15259 sky130_fd_sc_hd__dfbbn_1_2/a_891_329# V_LOW 2.26e-20
C15260 sky130_fd_sc_hd__nand2_8_3/A sky130_fd_sc_hd__nand2_8_3/Y 0.0776f
C15261 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# sky130_fd_sc_hd__inv_1_57/Y 0.0169f
C15262 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# sky130_fd_sc_hd__conb_1_49/HI 1.36e-20
C15263 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_1363_47# -2.65e-20
C15264 sky130_fd_sc_hd__dfbbn_1_37/a_1340_413# V_GND 2.04e-19
C15265 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0372f
C15266 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# V_GND 0.00331f
C15267 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.94e-19
C15268 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__inv_1_99/Y 1.64e-19
C15269 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# V_LOW 1.38e-19
C15270 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0398f
C15271 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0159f
C15272 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 5.11e-19
C15273 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# sky130_fd_sc_hd__inv_1_99/Y 5.43e-20
C15274 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# V_LOW 1.38e-19
C15275 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# V_GND -0.00543f
C15276 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__conb_1_24/LO 1.28e-20
C15277 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__conb_1_6/HI 0.00455f
C15278 FULL_COUNTER.COUNT_SUB_DFF8.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 6.91e-20
C15279 sky130_fd_sc_hd__inv_1_97/Y sky130_fd_sc_hd__inv_1_86/Y 0.0958f
C15280 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__conb_1_32/LO 8.09e-21
C15281 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__conb_1_0/HI 4.23e-19
C15282 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__conb_1_40/HI 0.02f
C15283 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0.00453f
C15284 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 5.15e-19
C15285 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 4.95e-19
C15286 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 2.4e-20
C15287 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.0109f
C15288 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 3.26e-20
C15289 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.366f
C15290 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__conb_1_9/HI 1.83e-19
C15291 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_50/a_791_47# 4.14e-20
C15292 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# -9.41e-19
C15293 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1672_329# -1.44e-20
C15294 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__inv_1_107/Y 1.03e-20
C15295 sky130_fd_sc_hd__dfbbn_1_22/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 7.09e-19
C15296 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# sky130_fd_sc_hd__conb_1_18/HI 3.29e-20
C15297 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.02e-19
C15298 sky130_fd_sc_hd__conb_1_36/HI sky130_fd_sc_hd__inv_1_108/Y 0.0018f
C15299 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# V_GND 0.00409f
C15300 sky130_fd_sc_hd__inv_1_5/Y V_LOW 0.13f
C15301 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF0.Q 2.14e-19
C15302 sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# V_GND 0.00103f
C15303 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__conb_1_38/HI 0.0133f
C15304 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# V_LOW -0.108f
C15305 sky130_fd_sc_hd__conb_1_5/HI sky130_fd_sc_hd__inv_16_2/Y 0.0011f
C15306 FALLING_COUNTER.COUNT_SUB_DFF14.Q FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0684f
C15307 sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# V_GND 9.97e-19
C15308 sky130_fd_sc_hd__conb_1_46/HI V_GND 0.137f
C15309 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0046f
C15310 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# V_LOW -0.109f
C15311 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 8.63e-20
C15312 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 7.25e-19
C15313 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__conb_1_39/LO 8.84e-20
C15314 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# -1.17e-19
C15315 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_20/Y 0.00357f
C15316 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_381_47# -0.00375f
C15317 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__inv_1_10/Y 1.8e-19
C15318 sky130_fd_sc_hd__inv_1_46/A V_LOW 0.471f
C15319 sky130_fd_sc_hd__inv_1_106/Y sky130_fd_sc_hd__conb_1_46/HI 0.0631f
C15320 sky130_fd_sc_hd__inv_1_79/A sky130_fd_sc_hd__inv_1_95/Y 0.00627f
C15321 RISING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_2/Y 1.35e-20
C15322 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 3.59e-22
C15323 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_39/A 1.76e-21
C15324 sky130_fd_sc_hd__dfbbn_1_26/a_1363_47# sky130_fd_sc_hd__conb_1_30/HI -4.88e-19
C15325 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 1.56e-21
C15326 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_64/A 0.0214f
C15327 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# sky130_fd_sc_hd__conb_1_51/HI 2.16e-20
C15328 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_381_47# -0.00419f
C15329 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# V_LOW -0.00147f
C15330 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 8.94e-21
C15331 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# V_GND -0.00489f
C15332 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF3.Q 1.44e-19
C15333 sky130_fd_sc_hd__dfbbn_1_25/a_1159_47# sky130_fd_sc_hd__conb_1_22/HI 4.8e-19
C15334 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# V_GND -0.00533f
C15335 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_40/A 0.185f
C15336 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_1_105/Y 0.0199f
C15337 sky130_fd_sc_hd__inv_1_45/A V_LOW 0.0768f
C15338 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.6e-20
C15339 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF5.Q 5.82e-20
C15340 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 9.16e-20
C15341 sky130_fd_sc_hd__dfbbn_1_10/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 8.36e-20
C15342 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_57/Y 0.0354f
C15343 sky130_fd_sc_hd__conb_1_24/HI sky130_fd_sc_hd__inv_1_58/Y 3.62e-20
C15344 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_581_47# 5.8e-19
C15345 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# sky130_fd_sc_hd__conb_1_12/HI -0.0126f
C15346 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_193_47# -0.0608f
C15347 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.00298f
C15348 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__conb_1_40/HI 0.018f
C15349 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 1.59e-19
C15350 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# V_LOW -9.94e-19
C15351 sky130_fd_sc_hd__inv_1_102/Y sky130_fd_sc_hd__conb_1_40/HI 0.102f
C15352 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# sky130_fd_sc_hd__inv_16_0/Y 4.34e-20
C15353 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1672_329# -1.44e-20
C15354 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0289f
C15355 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 1.29e-19
C15356 sky130_fd_sc_hd__dfbbn_1_0/a_891_329# V_GND 3.29e-19
C15357 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_22/Y 0.282f
C15358 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF0.Q 3.44e-20
C15359 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00284f
C15360 sky130_fd_sc_hd__inv_1_55/Y RISING_COUNTER.COUNT_SUB_DFF6.Q 2.94e-20
C15361 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF13.Q 4.21e-19
C15362 sky130_fd_sc_hd__inv_1_72/A sky130_fd_sc_hd__inv_1_76/A 0.191f
C15363 sky130_fd_sc_hd__inv_1_119/Y sky130_fd_sc_hd__inv_1_67/Y 4.56e-21
C15364 sky130_fd_sc_hd__dfbbn_1_50/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 8.97e-19
C15365 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# 0.00901f
C15366 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.0126f
C15367 sky130_fd_sc_hd__nand2_8_6/a_27_47# V_GND 0.0114f
C15368 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__conb_1_40/HI 1.9e-20
C15369 sky130_fd_sc_hd__dfbbn_1_7/a_891_329# sky130_fd_sc_hd__inv_1_18/Y 0.0036f
C15370 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00265f
C15371 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_18/HI 0.00148f
C15372 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0217f
C15373 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# V_GND 0.0046f
C15374 sky130_fd_sc_hd__inv_1_91/A Reset 0.0493f
C15375 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -7.6e-19
C15376 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# -0.00226f
C15377 sky130_fd_sc_hd__dfbbn_1_46/a_581_47# sky130_fd_sc_hd__inv_1_99/Y 2.34e-19
C15378 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00541f
C15379 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.42e-19
C15380 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__conb_1_32/HI 0.0104f
C15381 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# sky130_fd_sc_hd__conb_1_15/LO 8.84e-20
C15382 sky130_fd_sc_hd__dfbbn_1_33/a_1112_329# sky130_fd_sc_hd__conb_1_35/HI 0.00358f
C15383 sky130_fd_sc_hd__dfbbn_1_23/a_1363_47# V_GND 1.64e-19
C15384 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__inv_1_54/Y 8.18e-21
C15385 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 1.6e-20
C15386 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# -9.25e-19
C15387 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# -0.0103f
C15388 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# Reset 2.22e-19
C15389 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 1.3e-19
C15390 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 4.83e-21
C15391 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__nand2_8_4/a_27_47# 9.56e-19
C15392 sky130_fd_sc_hd__dfbbn_1_51/a_1672_329# sky130_fd_sc_hd__conb_1_40/HI 3.98e-19
C15393 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 2.27e-19
C15394 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__conb_1_27/LO 7.66e-19
C15395 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 3.84e-21
C15396 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 3.84e-21
C15397 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# sky130_fd_sc_hd__inv_1_107/Y 3.27e-19
C15398 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00776f
C15399 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.28e-20
C15400 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__inv_1_98/Y 6.01e-21
C15401 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 1.57e-19
C15402 sky130_fd_sc_hd__inv_1_110/Y V_GND 0.272f
C15403 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 2.53e-21
C15404 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__conb_1_1/HI 3.24e-19
C15405 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 2.59e-19
C15406 sky130_fd_sc_hd__inv_1_19/Y FULL_COUNTER.COUNT_SUB_DFF16.Q 1.56e-20
C15407 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.46e-20
C15408 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_4/Y 0.0769f
C15409 sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# V_LOW -2.68e-19
C15410 FALLING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_1/Y 0.17f
C15411 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# V_GND -0.0148f
C15412 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.67e-20
C15413 sky130_fd_sc_hd__dfbbn_1_47/a_1672_329# V_LOW -9.94e-19
C15414 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 1.07e-19
C15415 sky130_fd_sc_hd__inv_1_34/A V_SENSE 0.116f
C15416 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.43e-21
C15417 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00509f
C15418 sky130_fd_sc_hd__inv_1_93/A RISING_COUNTER.COUNT_SUB_DFF4.Q 0.00727f
C15419 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_16_2/Y 0.874f
C15420 sky130_fd_sc_hd__dfbbn_1_2/Q_N FULL_COUNTER.COUNT_SUB_DFF2.Q 9.2e-20
C15421 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# -0.00107f
C15422 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 5.59e-20
C15423 sky130_fd_sc_hd__nand3_1_0/a_109_47# V_LOW -2.94e-19
C15424 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 5.37e-22
C15425 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# -0.00138f
C15426 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -7.6e-19
C15427 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# -5.54e-21
C15428 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# sky130_fd_sc_hd__conb_1_17/HI 0.0204f
C15429 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# -1.44e-20
C15430 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# V_LOW -2.78e-35
C15431 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00104f
C15432 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# V_GND -3.6e-19
C15433 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 9.55e-21
C15434 sky130_fd_sc_hd__conb_1_5/LO V_GND -0.00203f
C15435 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0058f
C15436 sky130_fd_sc_hd__conb_1_27/LO sky130_fd_sc_hd__inv_16_0/Y 0.00673f
C15437 sky130_fd_sc_hd__dfbbn_1_47/a_1363_47# V_GND -3.72e-19
C15438 sky130_fd_sc_hd__conb_1_11/HI V_GND -0.201f
C15439 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# sky130_fd_sc_hd__inv_1_55/Y 0.00531f
C15440 sky130_fd_sc_hd__inv_1_66/Y CLOCK_GEN.SR_Op.Q 1.44e-19
C15441 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__nand3_1_0/Y 0.0782f
C15442 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.52e-20
C15443 sky130_fd_sc_hd__inv_1_64/Y V_LOW 0.0494f
C15444 sky130_fd_sc_hd__nand2_8_6/a_27_47# sky130_fd_sc_hd__nand3_1_1/Y 4.38e-19
C15445 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# V_LOW -0.115f
C15446 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0.0133f
C15447 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# V_LOW 0.00518f
C15448 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# sky130_fd_sc_hd__inv_1_12/Y 0.04f
C15449 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 1.5e-19
C15450 sky130_fd_sc_hd__inv_1_93/A sky130_fd_sc_hd__inv_1_65/Y 8.02e-20
C15451 sky130_fd_sc_hd__inv_1_70/A sky130_fd_sc_hd__inv_1_63/Y 1.32e-19
C15452 CLOCK_GEN.SR_Op.Q V_GND 1.15f
C15453 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1159_47# 0.00142f
C15454 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__inv_1_57/Y 0.226f
C15455 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 0.0201f
C15456 sky130_fd_sc_hd__inv_1_16/Y sky130_fd_sc_hd__conb_1_9/HI 4.52e-20
C15457 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0145f
C15458 sky130_fd_sc_hd__dfbbn_1_25/a_891_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00123f
C15459 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.00978f
C15460 sky130_fd_sc_hd__dfbbn_1_38/Q_N FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0192f
C15461 sky130_fd_sc_hd__nand2_8_8/a_27_47# sky130_fd_sc_hd__inv_1_66/Y 1.18e-20
C15462 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# 1.71e-20
C15463 sky130_fd_sc_hd__inv_1_72/Y V_LOW 0.108f
C15464 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_891_329# 3.9e-22
C15465 Reset sky130_fd_sc_hd__inv_16_1/Y 0.459f
C15466 sky130_fd_sc_hd__inv_1_95/A sky130_fd_sc_hd__inv_1_70/A 1.43e-19
C15467 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0022f
C15468 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.52e-21
C15469 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_1_100/Y 6.2e-21
C15470 sky130_fd_sc_hd__dfbbn_1_12/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.16e-19
C15471 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 0.0298f
C15472 sky130_fd_sc_hd__nand2_8_8/a_27_47# V_GND -0.00721f
C15473 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF15.Q 7.16e-19
C15474 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# V_GND 0.00157f
C15475 sky130_fd_sc_hd__dfbbn_1_41/a_891_329# V_GND 4.23e-19
C15476 sky130_fd_sc_hd__inv_1_75/A V_GND 0.92f
C15477 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# V_LOW 0.0073f
C15478 RISING_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__inv_1_61/Y 0.0172f
C15479 sky130_fd_sc_hd__dfbbn_1_1/a_891_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.1e-21
C15480 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# sky130_fd_sc_hd__inv_1_112/Y 2.65e-20
C15481 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0405f
C15482 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_1340_413# -6.8e-19
C15483 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__nand3_1_2/Y 0.382f
C15484 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__conb_1_2/LO 0.00107f
C15485 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_1_107/Y 0.00111f
C15486 sky130_fd_sc_hd__inv_1_51/A sky130_fd_sc_hd__nand2_8_1/a_27_47# 0.0202f
C15487 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0039f
C15488 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 1.27e-19
C15489 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# -5.33e-20
C15490 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_557_413# -3.67e-20
C15491 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# Reset 0.00256f
C15492 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# Reset 7.3e-19
C15493 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 0.00167f
C15494 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_43/LO 0.0374f
C15495 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_24/a_473_413# 4.79e-19
C15496 sky130_fd_sc_hd__conb_1_15/LO sky130_fd_sc_hd__inv_1_20/Y 1.19e-19
C15497 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# sky130_fd_sc_hd__inv_1_55/Y 0.00352f
C15498 sky130_fd_sc_hd__dfbbn_1_24/a_891_329# V_GND 3.37e-19
C15499 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00101f
C15500 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__conb_1_21/HI 0.00884f
C15501 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_5/LO 4.77e-20
C15502 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__conb_1_17/LO 0.00439f
C15503 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# sky130_fd_sc_hd__conb_1_11/HI 1.13e-21
C15504 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 0.00142f
C15505 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.42e-19
C15506 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# -2.33e-19
C15507 sky130_fd_sc_hd__conb_1_25/LO RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0176f
C15508 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# sky130_fd_sc_hd__inv_1_63/Y 1.56e-19
C15509 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -0.00592f
C15510 sky130_fd_sc_hd__inv_1_42/Y V_LOW 0.0962f
C15511 sky130_fd_sc_hd__conb_1_48/HI FALLING_COUNTER.COUNT_SUB_DFF10.Q 8.46e-19
C15512 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.83e-20
C15513 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# CLOCK_GEN.SR_Op.Q 2.71e-19
C15514 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# -9.32e-20
C15515 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0264f
C15516 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__conb_1_31/HI 0.171f
C15517 sky130_fd_sc_hd__dfbbn_1_12/a_1363_47# sky130_fd_sc_hd__conb_1_17/HI 4.96e-20
C15518 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.04e-19
C15519 sky130_fd_sc_hd__inv_1_56/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 4.64e-19
C15520 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand3_1_1/Y 4.33e-19
C15521 sky130_fd_sc_hd__dfbbn_1_0/Q_N V_LOW -0.00141f
C15522 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.87e-19
C15523 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0087f
C15524 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_35/HI 0.00479f
C15525 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_80/A 0.118f
C15526 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# V_LOW -0.103f
C15527 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_381_47# -0.00375f
C15528 sky130_fd_sc_hd__inv_1_83/Y Reset 0.0094f
C15529 sky130_fd_sc_hd__nand3_1_0/a_193_47# sky130_fd_sc_hd__inv_1_70/A 1.99e-20
C15530 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 0.00322f
C15531 sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# V_LOW -2.68e-19
C15532 sky130_fd_sc_hd__conb_1_46/LO sky130_fd_sc_hd__conb_1_46/HI 0.00393f
C15533 sky130_fd_sc_hd__dfbbn_1_47/a_1340_413# sky130_fd_sc_hd__inv_1_57/Y 1.9e-19
C15534 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_22/Y 1.69e-19
C15535 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.57e-20
C15536 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# sky130_fd_sc_hd__inv_16_1/Y 0.0354f
C15537 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 1.84e-19
C15538 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__inv_1_107/Y 0.117f
C15539 sky130_fd_sc_hd__dfbbn_1_45/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 2.14e-19
C15540 sky130_fd_sc_hd__dfbbn_1_18/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF7.Q 5.62e-19
C15541 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 6.25e-21
C15542 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0.00109f
C15543 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 2.88e-19
C15544 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 2.42e-19
C15545 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 1.08e-19
C15546 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 1.78e-21
C15547 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 1.78e-21
C15548 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 8.63e-20
C15549 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 0.00574f
C15550 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__inv_1_102/Y 1.49e-19
C15551 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 3.88e-20
C15552 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/Q_N 1.84e-19
C15553 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0.0122f
C15554 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 4.89e-21
C15555 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# V_LOW 0.0159f
C15556 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__conb_1_39/LO 0.015f
C15557 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__conb_1_4/HI 0.00621f
C15558 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# V_GND 0.00346f
C15559 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.00449f
C15560 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 8.79e-21
C15561 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 4.81e-21
C15562 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 6.25e-19
C15563 FULL_COUNTER.COUNT_SUB_DFF7.Q sky130_fd_sc_hd__conb_1_6/HI 6.56e-19
C15564 sky130_fd_sc_hd__dfbbn_1_33/a_1363_47# V_GND 1.64e-19
C15565 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0232f
C15566 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/Q_N -4.33e-20
C15567 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# V_LOW -2.78e-35
C15568 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# 3.86e-19
C15569 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# sky130_fd_sc_hd__inv_1_107/Y 0.00271f
C15570 sky130_fd_sc_hd__inv_1_91/A sky130_fd_sc_hd__inv_1_85/Y 0.07f
C15571 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__conb_1_7/LO 0.0116f
C15572 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# sky130_fd_sc_hd__nand3_1_2/Y 3.72e-19
C15573 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.1e-20
C15574 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__conb_1_31/HI 0.0177f
C15575 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# V_GND 2.54e-19
C15576 sky130_fd_sc_hd__conb_1_29/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 1.64e-20
C15577 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__conb_1_0/HI 2.87e-19
C15578 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__conb_1_1/HI 6.43e-19
C15579 sky130_fd_sc_hd__dfbbn_1_32/a_557_413# V_GND 2.69e-19
C15580 sky130_fd_sc_hd__dfbbn_1_11/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00268f
C15581 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 2.13e-19
C15582 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.58e-19
C15583 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_76/A 0.108f
C15584 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# sky130_fd_sc_hd__inv_1_103/Y 1.56e-20
C15585 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__conb_1_2/HI 6.43e-20
C15586 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_19/HI 0.0986f
C15587 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__conb_1_36/HI 0.0364f
C15588 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.00364f
C15589 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# Reset 3.79e-19
C15590 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 3.34e-20
C15591 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__inv_1_61/Y 3.09e-20
C15592 sky130_fd_sc_hd__dfbbn_1_22/a_557_413# sky130_fd_sc_hd__inv_1_61/Y 8.17e-19
C15593 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# sky130_fd_sc_hd__conb_1_11/HI 0.029f
C15594 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_97/Y 3.58e-20
C15595 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# sky130_fd_sc_hd__conb_1_34/HI 0.00306f
C15596 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_23/LO 0.0147f
C15597 FALLING_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_99/Y 0.0103f
C15598 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__conb_1_23/LO 8.81e-20
C15599 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00212f
C15600 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__conb_1_42/HI 0.0249f
C15601 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# sky130_fd_sc_hd__conb_1_45/HI 0.00166f
C15602 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__conb_1_38/HI 2.93e-19
C15603 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__conb_1_42/LO 8.09e-21
C15604 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF10.Q 9.32e-20
C15605 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__conb_1_32/HI 1.59e-19
C15606 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# sky130_fd_sc_hd__inv_1_59/Y 0.00195f
C15607 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI -5.14e-19
C15608 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0.0318f
C15609 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# RISING_COUNTER.COUNT_SUB_DFF9.Q 4.66e-19
C15610 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00604f
C15611 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.0246f
C15612 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# -1.66e-19
C15613 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_1672_329# -7.17e-20
C15614 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 0.0398f
C15615 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# sky130_fd_sc_hd__inv_1_103/Y 4.83e-20
C15616 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__conb_1_2/HI 6.13e-20
C15617 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# CLOCK_GEN.SR_Op.Q 2.03e-19
C15618 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# -3.72e-19
C15619 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# -0.00144f
C15620 sky130_fd_sc_hd__dfbbn_1_33/Q_N sky130_fd_sc_hd__conb_1_47/HI 2.18e-20
C15621 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.12e-22
C15622 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__inv_1_102/Y 0.00482f
C15623 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/Q_N -4.78e-20
C15624 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0499f
C15625 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 4.05e-19
C15626 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 0.19f
C15627 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 0.00298f
C15628 sky130_fd_sc_hd__dfbbn_1_35/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 4.74e-19
C15629 sky130_fd_sc_hd__conb_1_40/LO sky130_fd_sc_hd__conb_1_51/HI 0.0156f
C15630 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__inv_1_108/Y 0.00145f
C15631 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# sky130_fd_sc_hd__inv_1_4/Y 1.07e-20
C15632 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 2.22e-20
C15633 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 0.0025f
C15634 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 7.65e-21
C15635 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# sky130_fd_sc_hd__conb_1_27/HI 3.9e-19
C15636 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# V_LOW -2.68e-19
C15637 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 4.65e-21
C15638 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 7.87e-20
C15639 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 0.00384f
C15640 sky130_fd_sc_hd__inv_1_97/Y V_GND 0.129f
C15641 sky130_fd_sc_hd__dfbbn_1_48/a_891_329# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00109f
C15642 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.22e-20
C15643 sky130_fd_sc_hd__dfbbn_1_41/Q_N V_LOW -0.00245f
C15644 sky130_fd_sc_hd__inv_1_107/Y sky130_fd_sc_hd__inv_16_0/Y 4.78e-21
C15645 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 0.00188f
C15646 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 3.74e-20
C15647 sky130_fd_sc_hd__nand2_8_3/Y sky130_fd_sc_hd__inv_1_75/A 0.0963f
C15648 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_16_2/Y 0.95f
C15649 FULL_COUNTER.COUNT_SUB_DFF16.Q sky130_fd_sc_hd__conb_1_12/HI 0.174f
C15650 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 7.28e-21
C15651 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_9/a_791_47# 6.08e-19
C15652 sky130_fd_sc_hd__dfbbn_1_10/a_1112_329# V_LOW -0.00266f
C15653 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_64/A 3.78e-19
C15654 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_1_11/Y 3.86e-20
C15655 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# V_LOW 0.0101f
C15656 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 3.04e-19
C15657 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 1.15e-20
C15658 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 3.64e-20
C15659 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__conb_1_42/HI 0.00802f
C15660 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__conb_1_30/HI 5.77e-21
C15661 sky130_fd_sc_hd__dfbbn_1_16/a_1159_47# sky130_fd_sc_hd__conb_1_4/HI 2.09e-19
C15662 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 3.16e-19
C15663 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# sky130_fd_sc_hd__dfbbn_1_3/a_791_47# 2.69e-19
C15664 sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# V_GND 2.83e-19
C15665 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0444f
C15666 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_16_1/Y 0.00102f
C15667 sky130_fd_sc_hd__conb_1_24/LO CLOCK_GEN.SR_Op.Q 3.4e-21
C15668 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# sky130_fd_sc_hd__inv_1_58/Y 2.37e-19
C15669 sky130_fd_sc_hd__dfbbn_1_27/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00119f
C15670 sky130_fd_sc_hd__nand2_8_9/Y V_LOW 0.0781f
C15671 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__conb_1_38/HI 8.33e-19
C15672 sky130_fd_sc_hd__dfbbn_1_24/Q_N V_LOW -2.68e-19
C15673 FALLING_COUNTER.COUNT_SUB_DFF1.Q FALLING_COUNTER.COUNT_SUB_DFF0.Q 1.62f
C15674 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 0.221f
C15675 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0418f
C15676 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_16_0/Y 0.291f
C15677 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_10/HI 0.00276f
C15678 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0189f
C15679 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# 0.00147f
C15680 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# V_LOW -0.318f
C15681 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# sky130_fd_sc_hd__conb_1_31/HI 0.00242f
C15682 sky130_fd_sc_hd__dfbbn_1_10/a_581_47# V_GND -9.18e-19
C15683 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# -3.07e-19
C15684 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# -2.32e-19
C15685 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# sky130_fd_sc_hd__conb_1_36/HI 0.00333f
C15686 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# sky130_fd_sc_hd__conb_1_1/HI -0.0112f
C15687 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__inv_1_66/Y 0.0792f
C15688 RISING_COUNTER.COUNT_SUB_DFF12.Q CLOCK_GEN.SR_Op.Q 0.00403f
C15689 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 9.4e-21
C15690 sky130_fd_sc_hd__dfbbn_1_40/a_1672_329# sky130_fd_sc_hd__conb_1_36/HI 9.52e-19
C15691 FALLING_COUNTER.COUNT_SUB_DFF1.Q V_LOW 1.24f
C15692 RISING_COUNTER.COUNT_SUB_DFF11.Q sky130_fd_sc_hd__conb_1_22/HI 0.00149f
C15693 RISING_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_53/Y 1.31e-20
C15694 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_22/Y 3.42e-20
C15695 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_22/a_647_21# 1.75e-19
C15696 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 3.42e-19
C15697 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# sky130_fd_sc_hd__inv_1_5/Y 1.43e-19
C15698 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.125f
C15699 sky130_fd_sc_hd__inv_1_96/Y V_GND 0.07f
C15700 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# V_LOW 0.0173f
C15701 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# V_GND 0.00776f
C15702 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# V_LOW 0.067f
C15703 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 0.0025f
C15704 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# V_GND -0.0442f
C15705 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__conb_1_13/HI 0.00964f
C15706 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# sky130_fd_sc_hd__inv_1_10/Y 0.00665f
C15707 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__conb_1_40/HI 9.3e-19
C15708 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# sky130_fd_sc_hd__conb_1_24/HI 9.37e-21
C15709 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 0.0578f
C15710 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 8.64e-21
C15711 sky130_fd_sc_hd__dfbbn_1_46/a_1159_47# sky130_fd_sc_hd__inv_16_1/Y 0.00472f
C15712 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# sky130_fd_sc_hd__inv_1_103/Y 7.15e-19
C15713 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_1672_329# -5.16e-20
C15714 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# -1.66e-19
C15715 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.0298f
C15716 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_91/Y 1.2e-19
C15717 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 1.86e-21
C15718 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.01e-20
C15719 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00191f
C15720 sky130_fd_sc_hd__inv_1_69/Y V_GND 0.614f
C15721 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# V_GND 0.00774f
C15722 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.29e-21
C15723 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# V_GND 0.0111f
C15724 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00185f
C15725 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# V_GND -0.00166f
C15726 sky130_fd_sc_hd__inv_1_68/Y V_GND 0.00474f
C15727 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_112/Y 5.79e-20
C15728 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# sky130_fd_sc_hd__inv_1_21/Y 0.00253f
C15729 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.514f
C15730 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 9.22e-20
C15731 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 9.07e-21
C15732 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# sky130_fd_sc_hd__conb_1_27/HI 2.99e-19
C15733 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 9.12e-19
C15734 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# V_LOW -0.323f
C15735 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 1.81e-20
C15736 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_107/Y 1.68e-20
C15737 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.0194f
C15738 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00175f
C15739 sky130_fd_sc_hd__inv_1_85/Y sky130_fd_sc_hd__inv_1_83/Y 0.118f
C15740 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.29e-19
C15741 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# -1.98e-19
C15742 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# -2.52e-19
C15743 Reset V_LOW 2.54f
C15744 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 1.06e-19
C15745 sky130_fd_sc_hd__inv_1_51/Y V_GND -0.00301f
C15746 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 8.78e-21
C15747 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0.003f
C15748 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 6.66e-19
C15749 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 8.4e-21
C15750 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 9.05e-19
C15751 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 9.75e-20
C15752 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__conb_1_22/HI 0.00233f
C15753 sky130_fd_sc_hd__dfbbn_1_32/Q_N FALLING_COUNTER.COUNT_SUB_DFF6.Q 5.44e-20
C15754 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_76/A 4.73e-19
C15755 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__conb_1_16/LO 0.00366f
C15756 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_19/a_891_329# 1.93e-21
C15757 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 1.85f
C15758 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# V_GND -0.0486f
C15759 sky130_fd_sc_hd__dfbbn_1_34/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF12.Q 0.00174f
C15760 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# sky130_fd_sc_hd__inv_2_0/Y 3.77e-20
C15761 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_34/a_557_413# -0.0012f
C15762 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# -0.0244f
C15763 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# sky130_fd_sc_hd__inv_1_58/Y 4.07e-20
C15764 sky130_fd_sc_hd__conb_1_7/HI FULL_COUNTER.COUNT_SUB_DFF8.Q 0.0763f
C15765 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.00286f
C15766 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_16_0/Y 0.0187f
C15767 sky130_fd_sc_hd__dfbbn_1_48/a_1112_329# V_LOW 4.8e-20
C15768 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.55e-21
C15769 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# V_LOW -0.0995f
C15770 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# sky130_fd_sc_hd__conb_1_27/HI 8.55e-20
C15771 sky130_fd_sc_hd__dfbbn_1_39/Q_N sky130_fd_sc_hd__inv_1_107/Y 5.93e-20
C15772 sky130_fd_sc_hd__inv_1_96/Y sky130_fd_sc_hd__nand3_1_1/Y 7.33e-19
C15773 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# 0.00243f
C15774 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.0417f
C15775 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# sky130_fd_sc_hd__inv_16_0/Y 7.37e-19
C15776 sky130_fd_sc_hd__inv_1_7/Y V_LOW 0.0955f
C15777 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.22e-20
C15778 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# V_LOW -1.21e-19
C15779 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00684f
C15780 RISING_COUNTER.COUNT_SUB_DFF3.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0245f
C15781 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 8e-21
C15782 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0.00819f
C15783 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_13/Y 1.59e-20
C15784 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# -7.17e-20
C15785 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# -1.64e-19
C15786 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__conb_1_19/LO 4.01e-19
C15787 sky130_fd_sc_hd__dfbbn_1_37/Q_N sky130_fd_sc_hd__inv_1_103/Y 2.81e-21
C15788 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 6.47e-19
C15789 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# V_LOW -0.317f
C15790 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# sky130_fd_sc_hd__conb_1_47/HI 7.46e-20
C15791 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_51/a_891_329# 2.22e-21
C15792 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.34e-19
C15793 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# sky130_fd_sc_hd__inv_1_5/Y 3.01e-19
C15794 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1_26/Y 0.0421f
C15795 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_31/A 0.103f
C15796 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_1/Y 0.178f
C15797 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0632f
C15798 sky130_fd_sc_hd__conb_1_11/LO V_LOW 0.0645f
C15799 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__inv_16_2/Y 0.0144f
C15800 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 0.00214f
C15801 sky130_fd_sc_hd__dfbbn_1_48/a_581_47# V_GND 1.58e-19
C15802 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# -0.0242f
C15803 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__dfbbn_1_29/a_557_413# -3.67e-20
C15804 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# V_LOW -0.00121f
C15805 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# V_GND 0.00178f
C15806 sky130_fd_sc_hd__nand2_1_0/a_113_47# V_GND -8.04e-20
C15807 sky130_fd_sc_hd__dfbbn_1_8/a_1340_413# V_LOW 2.94e-20
C15808 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__dfbbn_1_11/a_473_413# -0.00312f
C15809 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_647_21# -0.00746f
C15810 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 0.002f
C15811 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 2.11e-21
C15812 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 2.73e-21
C15813 sky130_fd_sc_hd__dfbbn_1_12/a_891_329# V_GND 3.13e-19
C15814 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 0.0235f
C15815 sky130_fd_sc_hd__dfbbn_1_34/a_1672_329# V_GND 1.58e-19
C15816 sky130_fd_sc_hd__conb_1_12/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0469f
C15817 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# -6.23e-21
C15818 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_8/a_381_47# -0.00832f
C15819 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.00233f
C15820 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# V_LOW 0.0125f
C15821 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__dfbbn_1_39/a_193_47# -0.141f
C15822 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__conb_1_37/HI 6.22e-20
C15823 sky130_fd_sc_hd__dfbbn_1_22/Q_N RISING_COUNTER.COUNT_SUB_DFF9.Q 0.00306f
C15824 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# V_GND 0.00781f
C15825 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 1.02e-19
C15826 sky130_fd_sc_hd__inv_1_40/A V_GND 0.0819f
C15827 sky130_fd_sc_hd__inv_1_67/Y sky130_fd_sc_hd__nand2_1_0/Y 1.76e-19
C15828 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_62/Y 1.31e-19
C15829 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 4.86e-19
C15830 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 3.66e-19
C15831 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# -0.0071f
C15832 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.014f
C15833 sky130_fd_sc_hd__dfbbn_1_42/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF7.Q 6.03e-20
C15834 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__conb_1_27/HI 5.7e-20
C15835 sky130_fd_sc_hd__dfbbn_1_29/a_1672_329# V_GND 3.58e-19
C15836 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# V_GND 0.00387f
C15837 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# V_LOW 0.0204f
C15838 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.08e-20
C15839 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# V_LOW 0.00685f
C15840 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# sky130_fd_sc_hd__conb_1_44/HI 0.00692f
C15841 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_27_47# 0.0346f
C15842 sky130_fd_sc_hd__dfbbn_1_8/a_1159_47# V_GND -0.0016f
C15843 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__conb_1_36/LO 0.00107f
C15844 FULL_COUNTER.COUNT_SUB_DFF6.Q V_LOW 3.15f
C15845 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# V_LOW -0.00288f
C15846 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_78/A 0.026f
C15847 sky130_fd_sc_hd__dfbbn_1_17/Q_N sky130_fd_sc_hd__inv_1_4/Y 5.85e-22
C15848 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0322f
C15849 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 3.82e-19
C15850 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_15/a_581_47# 2.86e-19
C15851 sky130_fd_sc_hd__dfbbn_1_40/a_557_413# V_GND 3.32e-19
C15852 sky130_fd_sc_hd__inv_1_57/Y V_LOW 0.136f
C15853 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 4.32e-20
C15854 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00101f
C15855 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# sky130_fd_sc_hd__conb_1_23/LO 3.81e-20
C15856 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.0138f
C15857 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 6.01e-19
C15858 sky130_fd_sc_hd__conb_1_25/LO sky130_fd_sc_hd__conb_1_26/LO 0.00434f
C15859 sky130_fd_sc_hd__inv_1_14/Y sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 4.44e-20
C15860 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# -1.76e-19
C15861 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# sky130_fd_sc_hd__dfbbn_1_20/a_941_21# -0.0137f
C15862 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# sky130_fd_sc_hd__dfbbn_1_20/a_473_413# -0.012f
C15863 sky130_fd_sc_hd__dfbbn_1_29/a_557_413# Reset 8.26e-19
C15864 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 4.11e-21
C15865 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_22/HI 0.277f
C15866 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# V_GND 1.81e-19
C15867 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# sky130_fd_sc_hd__inv_1_21/Y 1.05e-19
C15868 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 0.0161f
C15869 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# sky130_fd_sc_hd__conb_1_22/HI 0.00191f
C15870 sky130_fd_sc_hd__dfbbn_1_16/a_891_329# V_GND 4.66e-19
C15871 sky130_fd_sc_hd__dfbbn_1_38/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF9.Q 8.52e-19
C15872 RISING_COUNTER.COUNT_SUB_DFF13.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 1.02f
C15873 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__conb_1_51/LO 0.134f
C15874 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# sky130_fd_sc_hd__dfbbn_1_12/a_381_47# -0.00516f
C15875 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# V_GND 2.98e-19
C15876 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_56/Y 3.03e-19
C15877 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.0138f
C15878 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# V_LOW -0.00447f
C15879 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.69e-19
C15880 sky130_fd_sc_hd__dfbbn_1_36/a_1672_329# V_GND 1.7e-19
C15881 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_25/LO 4.54e-20
C15882 sky130_fd_sc_hd__dfbbn_1_42/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.53e-19
C15883 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0518f
C15884 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_19/Y 2.62e-20
C15885 sky130_fd_sc_hd__dfbbn_1_20/a_1672_329# V_LOW -2.68e-19
C15886 sky130_fd_sc_hd__inv_1_70/Y sky130_fd_sc_hd__nand3_1_0/Y 0.077f
C15887 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 0.0151f
C15888 sky130_fd_sc_hd__dfbbn_1_41/a_1363_47# sky130_fd_sc_hd__conb_1_27/HI 4.22e-19
C15889 sky130_fd_sc_hd__dfbbn_1_22/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.00954f
C15890 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# sky130_fd_sc_hd__inv_1_21/Y 1.57e-20
C15891 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# sky130_fd_sc_hd__dfbbn_1_36/a_891_329# -1.42e-19
C15892 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# -0.0244f
C15893 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_557_413# -0.0012f
C15894 sky130_fd_sc_hd__dfbbn_1_3/Q_N FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00159f
C15895 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.0113f
C15896 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__conb_1_44/HI 0.0518f
C15897 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 4.87e-21
C15898 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# sky130_fd_sc_hd__conb_1_47/HI 0.0273f
C15899 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 2.76e-20
C15900 sky130_fd_sc_hd__dfbbn_1_40/a_1363_47# sky130_fd_sc_hd__conb_1_47/HI 1.2e-19
C15901 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# V_LOW 1.38e-19
C15902 sky130_fd_sc_hd__dfbbn_1_4/a_557_413# V_GND 1.65e-19
C15903 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# 0.00475f
C15904 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00135f
C15905 sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 6.19e-20
C15906 sky130_fd_sc_hd__dfbbn_1_6/a_557_413# sky130_fd_sc_hd__inv_1_12/Y 4.19e-20
C15907 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 4.68e-21
C15908 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# sky130_fd_sc_hd__inv_1_65/Y 0.00656f
C15909 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 4.86e-20
C15910 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 2.53e-19
C15911 sky130_fd_sc_hd__conb_1_31/HI RISING_COUNTER.COUNT_SUB_DFF5.Q 2.18e-19
C15912 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# -1.31e-19
C15913 sky130_fd_sc_hd__dfbbn_1_14/a_891_329# sky130_fd_sc_hd__inv_1_12/Y 2.92e-19
C15914 sky130_fd_sc_hd__dfbbn_1_20/a_1363_47# V_GND 1.88e-19
C15915 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# sky130_fd_sc_hd__conb_1_24/HI 9.64e-22
C15916 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 0.0252f
C15917 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 0.00497f
C15918 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__conb_1_43/LO 0.0627f
C15919 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 2.96e-21
C15920 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0.0175f
C15921 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00685f
C15922 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_28/a_1363_47# 7.69e-20
C15923 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# V_LOW 0.00666f
C15924 sky130_fd_sc_hd__inv_1_76/A V_SENSE 1.4f
C15925 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0165f
C15926 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# V_LOW -0.00223f
C15927 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# sky130_fd_sc_hd__conb_1_37/HI 1.33e-19
C15928 sky130_fd_sc_hd__inv_1_62/Y sky130_fd_sc_hd__conb_1_32/HI 0.0049f
C15929 sky130_fd_sc_hd__inv_1_52/Y RISING_COUNTER.COUNT_SUB_DFF2.Q 0.323f
C15930 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# sky130_fd_sc_hd__conb_1_32/HI 0.00733f
C15931 sky130_fd_sc_hd__dfbbn_1_1/a_1672_329# V_GND 2.24e-19
C15932 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF18.Q 5.45e-19
C15933 sky130_fd_sc_hd__inv_1_17/Y sky130_fd_sc_hd__conb_1_25/HI 1.36e-20
C15934 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# V_LOW 0.0219f
C15935 sky130_fd_sc_hd__dfbbn_1_9/a_1112_329# V_GND 7.01e-19
C15936 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__inv_16_1/Y 4.47e-19
C15937 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__inv_16_0/Y 4.06e-21
C15938 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# 4.62e-19
C15939 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 1.15e-19
C15940 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# 6.21e-20
C15941 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 6.15e-20
C15942 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 2.35e-19
C15943 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# RISING_COUNTER.COUNT_SUB_DFF10.Q 5.01e-19
C15944 FULL_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__inv_1_9/Y 0.177f
C15945 FALLING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_39/LO 0.0142f
C15946 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# sky130_fd_sc_hd__dfbbn_1_40/a_941_21# -1.42e-32
C15947 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# -1.85e-19
C15948 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# -5.54e-21
C15949 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__inv_1_71/A 0.0174f
C15950 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.19e-21
C15951 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# V_LOW -1.39e-35
C15952 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# 3.78e-19
C15953 sky130_fd_sc_hd__dfbbn_1_34/a_1159_47# sky130_fd_sc_hd__conb_1_44/HI -0.00262f
C15954 sky130_fd_sc_hd__dfbbn_1_23/Q_N RISING_COUNTER.COUNT_SUB_DFF7.Q 0.00109f
C15955 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.077f
C15956 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# V_GND 0.0557f
C15957 FULL_COUNTER.COUNT_SUB_DFF12.Q FULL_COUNTER.COUNT_SUB_DFF4.Q 0.846f
C15958 sky130_fd_sc_hd__conb_1_14/HI V_LOW 0.171f
C15959 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# V_LOW -1.39e-35
C15960 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 4.45e-20
C15961 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# V_GND -0.00464f
C15962 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 1.49e-19
C15963 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_2/HI 0.0258f
C15964 sky130_fd_sc_hd__inv_1_103/Y sky130_fd_sc_hd__inv_1_105/Y 9.26e-22
C15965 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_50/A 0.0696f
C15966 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 3.65e-21
C15967 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 2.71e-19
C15968 sky130_fd_sc_hd__inv_1_68/A V_LOW 0.513f
C15969 sky130_fd_sc_hd__dfbbn_1_25/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.0266f
C15970 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 5.14e-19
C15971 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0.00112f
C15972 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 1.16e-19
C15973 sky130_fd_sc_hd__dfbbn_1_49/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0257f
C15974 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# sky130_fd_sc_hd__conb_1_41/HI 1.25e-21
C15975 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 1.1e-19
C15976 sky130_fd_sc_hd__dfbbn_1_7/a_557_413# V_GND 1.37e-19
C15977 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__conb_1_18/LO 1.29e-19
C15978 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__conb_1_45/HI 1.1e-19
C15979 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 0.00636f
C15980 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_647_21# -0.00108f
C15981 sky130_fd_sc_hd__conb_1_1/LO sky130_fd_sc_hd__inv_16_2/Y 0.00103f
C15982 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# -9.41e-19
C15983 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00996f
C15984 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 3.58e-19
C15985 sky130_fd_sc_hd__inv_1_85/Y V_LOW 0.14f
C15986 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 7.28e-19
C15987 sky130_fd_sc_hd__conb_1_4/HI sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 6.53e-20
C15988 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# -0.00107f
C15989 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# -1.6e-19
C15990 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# -5.54e-21
C15991 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_1_98/Y 1.1e-19
C15992 sky130_fd_sc_hd__conb_1_8/LO V_LOW 0.0879f
C15993 sky130_fd_sc_hd__inv_1_104/Y FALLING_COUNTER.COUNT_SUB_DFF11.Q 8.9e-19
C15994 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 0.0295f
C15995 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_16/a_381_47# -2.53e-20
C15996 sky130_fd_sc_hd__dfbbn_1_7/a_581_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00175f
C15997 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 0.0166f
C15998 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# V_LOW 0.00328f
C15999 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 8.63e-20
C16000 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 2.88e-19
C16001 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 1.08e-19
C16002 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 0.00109f
C16003 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 2.42e-19
C16004 sky130_fd_sc_hd__conb_1_3/LO V_GND 0.00376f
C16005 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 0.0301f
C16006 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_12/Y 0.133f
C16007 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.0024f
C16008 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# sky130_fd_sc_hd__dfbbn_1_14/a_381_47# -0.00869f
C16009 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF10.Q 3.09e-19
C16010 sky130_fd_sc_hd__conb_1_37/LO sky130_fd_sc_hd__inv_1_91/Y 1.87e-21
C16011 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__inv_1_10/Y 3.17e-20
C16012 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 4.95e-19
C16013 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 2.2e-19
C16014 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__inv_16_0/Y 0.125f
C16015 sky130_fd_sc_hd__dfbbn_1_12/Q_N V_LOW -0.0104f
C16016 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 2.12e-21
C16017 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# -0.00335f
C16018 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_1/a_557_413# -0.0012f
C16019 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 6.71e-19
C16020 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 4.56e-21
C16021 sky130_fd_sc_hd__dfbbn_1_27/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00169f
C16022 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.8e-19
C16023 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 1.8e-19
C16024 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0111f
C16025 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0.0111f
C16026 sky130_fd_sc_hd__inv_1_88/Y sky130_fd_sc_hd__dfbbn_1_48/a_891_329# 7.97e-21
C16027 sky130_fd_sc_hd__conb_1_27/LO V_GND -0.00238f
C16028 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.598f
C16029 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 6.77e-20
C16030 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 1.76e-20
C16031 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 3.34e-19
C16032 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 1.14e-19
C16033 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 1.8e-19
C16034 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# sky130_fd_sc_hd__inv_1_102/Y 4.19e-19
C16035 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# sky130_fd_sc_hd__conb_1_47/HI 0.0691f
C16036 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__inv_1_15/Y 1.45e-19
C16037 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# sky130_fd_sc_hd__conb_1_36/HI 3.05e-19
C16038 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# -1.56e-19
C16039 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.03e-23
C16040 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# sky130_fd_sc_hd__conb_1_22/HI 1.86e-20
C16041 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__dfbbn_1_11/a_381_47# 6.21e-21
C16042 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# sky130_fd_sc_hd__inv_16_0/Y 0.0113f
C16043 sky130_fd_sc_hd__conb_1_38/LO V_GND 0.0183f
C16044 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 0.0259f
C16045 sky130_fd_sc_hd__conb_1_50/LO sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 6.78e-21
C16046 FULL_COUNTER.COUNT_SUB_DFF1.Q FULL_COUNTER.COUNT_SUB_DFF13.Q 0.00528f
C16047 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 1.47e-21
C16048 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_35/a_1672_329# 1.09e-20
C16049 sky130_fd_sc_hd__inv_1_109/Y sky130_fd_sc_hd__conb_1_47/HI 1.03e-19
C16050 sky130_fd_sc_hd__dfbbn_1_13/a_557_413# V_LOW -9.15e-19
C16051 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_76/A 5.91e-19
C16052 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# 2.79e-19
C16053 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# V_GND -3.72e-21
C16054 sky130_fd_sc_hd__dfbbn_1_40/Q_N FALLING_COUNTER.COUNT_SUB_DFF6.Q 0.0212f
C16055 sky130_fd_sc_hd__dfbbn_1_31/Q_N sky130_fd_sc_hd__conb_1_37/HI 5.06e-19
C16056 FULL_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__inv_16_2/Y 1.37f
C16057 sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# sky130_fd_sc_hd__conb_1_32/HI 1.09e-20
C16058 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 1.06e-20
C16059 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_6/Y 0.00159f
C16060 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0362f
C16061 sky130_fd_sc_hd__inv_1_74/Y sky130_fd_sc_hd__inv_1_95/Y 8e-20
C16062 sky130_fd_sc_hd__conb_1_36/HI FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.83e-19
C16063 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# V_LOW 0.00353f
C16064 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# sky130_fd_sc_hd__inv_1_15/Y 5.37e-19
C16065 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__conb_1_2/LO 7.31e-20
C16066 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# 3.66e-22
C16067 sky130_fd_sc_hd__inv_1_56/Y V_LOW 0.102f
C16068 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# V_GND 0.014f
C16069 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 4.93e-20
C16070 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 4.93e-20
C16071 sky130_fd_sc_hd__conb_1_19/HI sky130_fd_sc_hd__dfbbn_1_17/Q_N 7.43e-21
C16072 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__inv_1_15/Y 0.00816f
C16073 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# -7.47e-20
C16074 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_1_60/Y 2.08e-19
C16075 sky130_fd_sc_hd__dfbbn_1_10/a_891_329# sky130_fd_sc_hd__inv_16_2/Y 2.78e-20
C16076 FALLING_COUNTER.COUNT_SUB_DFF4.Q sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 1.47e-21
C16077 sky130_fd_sc_hd__conb_1_8/HI V_GND -0.207f
C16078 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 8.91e-20
C16079 sky130_fd_sc_hd__dfbbn_1_16/Q_N V_LOW -0.0104f
C16080 sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00357f
C16081 sky130_fd_sc_hd__dfbbn_1_13/a_1340_413# V_GND 1.8e-19
C16082 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__inv_1_108/Y 0.0704f
C16083 sky130_fd_sc_hd__dfbbn_1_14/Q_N V_LOW -0.0104f
C16084 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# -2.01e-20
C16085 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# -7.6e-19
C16086 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# V_LOW 0.00676f
C16087 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# V_GND -0.00536f
C16088 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 0.0016f
C16089 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 8.59e-19
C16090 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF2.Q 2.67e-19
C16091 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 0.0577f
C16092 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00153f
C16093 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.87e-20
C16094 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__dfbbn_1_21/a_581_47# -2.6e-20
C16095 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 0.00111f
C16096 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__conb_1_48/LO 1.03e-19
C16097 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__inv_16_1/Y 1.09e-19
C16098 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__conb_1_18/LO 0.012f
C16099 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 7.44e-21
C16100 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 4.58e-19
C16101 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 2.38e-20
C16102 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 0.00127f
C16103 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 1.25e-19
C16104 sky130_fd_sc_hd__inv_1_17/Y FULL_COUNTER.COUNT_SUB_DFF3.Q 1.47e-19
C16105 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_71/A 1.49e-19
C16106 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF13.Q 5.26e-20
C16107 sky130_fd_sc_hd__dfbbn_1_49/a_891_329# V_GND 4.69e-19
C16108 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 3.15e-20
C16109 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# sky130_fd_sc_hd__conb_1_51/HI 3.13e-19
C16110 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_16/a_1672_329# -0.00148f
C16111 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_20/Y 8.62e-19
C16112 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 6.45e-19
C16113 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 2.48e-20
C16114 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 4.12e-19
C16115 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 1.62e-19
C16116 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 7.9e-19
C16117 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 2.27e-19
C16118 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__conb_1_50/HI 4.56e-21
C16119 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# V_LOW 0.00666f
C16120 sky130_fd_sc_hd__dfbbn_1_44/Q_N RISING_COUNTER.COUNT_SUB_DFF11.Q 1.01e-21
C16121 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 1.66e-20
C16122 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.66e-20
C16123 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# RISING_COUNTER.COUNT_SUB_DFF5.Q 8.85e-20
C16124 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_25/a_891_329# 1.3e-20
C16125 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__conb_1_33/LO 0.00178f
C16126 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 3.5e-19
C16127 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_647_21# 1.88e-21
C16128 sky130_fd_sc_hd__dfbbn_1_21/Q_N RISING_COUNTER.COUNT_SUB_DFF2.Q 2.47e-19
C16129 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# -0.00107f
C16130 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__conb_1_23/HI 1.27e-19
C16131 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0786f
C16132 sky130_fd_sc_hd__inv_1_20/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0013f
C16133 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 1.04e-20
C16134 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 1.04e-19
C16135 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00312f
C16136 sky130_fd_sc_hd__dfbbn_1_11/Q_N sky130_fd_sc_hd__inv_1_21/Y 1.26e-20
C16137 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 0.00124f
C16138 sky130_fd_sc_hd__dfbbn_1_5/a_1112_329# V_LOW -0.00266f
C16139 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 9.55e-22
C16140 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 9.55e-22
C16141 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# sky130_fd_sc_hd__dfbbn_1_9/a_891_329# -2.2e-20
C16142 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# -4.1e-19
C16143 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 6.77e-21
C16144 sky130_fd_sc_hd__inv_1_98/Y FALLING_COUNTER.COUNT_SUB_DFF8.Q 3.2e-21
C16145 sky130_fd_sc_hd__conb_1_33/LO RISING_COUNTER.COUNT_SUB_DFF0.Q 0.153f
C16146 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# V_LOW 1.38e-19
C16147 sky130_fd_sc_hd__dfbbn_1_5/a_891_329# sky130_fd_sc_hd__inv_1_13/Y 2.32e-20
C16148 sky130_fd_sc_hd__nand2_8_2/A sky130_fd_sc_hd__inv_1_78/A 0.00567f
C16149 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_10/Q_N 0.0014f
C16150 sky130_fd_sc_hd__dfbbn_1_16/a_557_413# sky130_fd_sc_hd__inv_1_8/Y 8.17e-19
C16151 sky130_fd_sc_hd__dfbbn_1_3/a_891_329# V_LOW 2.26e-20
C16152 sky130_fd_sc_hd__dfbbn_1_17/a_891_329# V_GND 4.11e-19
C16153 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_4/a_791_47# 0.00417f
C16154 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00313f
C16155 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_2/a_27_47# 0.0461f
C16156 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# sky130_fd_sc_hd__inv_1_76/A 1.87e-19
C16157 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.15e-19
C16158 sky130_fd_sc_hd__dfbbn_1_20/a_1112_329# sky130_fd_sc_hd__inv_1_53/Y 6.2e-19
C16159 sky130_fd_sc_hd__dfbbn_1_5/a_581_47# V_GND -9.06e-19
C16160 sky130_fd_sc_hd__conb_1_30/HI V_LOW 0.0414f
C16161 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 3.78e-19
C16162 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 7.87e-19
C16163 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 1.53e-19
C16164 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0.00187f
C16165 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 0.00247f
C16166 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 1.67e-19
C16167 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 7.63e-19
C16168 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.0405f
C16169 sky130_fd_sc_hd__dfbbn_1_11/Q_N FULL_COUNTER.COUNT_SUB_DFF18.Q 0.00135f
C16170 sky130_fd_sc_hd__inv_1_31/Y V_GND 0.0233f
C16171 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0328f
C16172 sky130_fd_sc_hd__dfbbn_1_43/a_1112_329# V_GND 8.21e-19
C16173 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 1.62e-20
C16174 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_647_21# -0.00618f
C16175 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# V_GND 0.00362f
C16176 sky130_fd_sc_hd__dfbbn_1_14/a_1672_329# sky130_fd_sc_hd__inv_1_15/Y 6.09e-21
C16177 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_40/Q_N -4.24e-20
C16178 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# RISING_COUNTER.COUNT_SUB_DFF3.Q 9.7e-21
C16179 sky130_fd_sc_hd__nand2_8_5/a_27_47# sky130_fd_sc_hd__nand3_1_0/a_193_47# 6.69e-20
C16180 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 2.79e-19
C16181 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# sky130_fd_sc_hd__inv_1_16/Y 2.55e-21
C16182 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_50/A 3.1e-19
C16183 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__inv_1_16/Y 0.00248f
C16184 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# -2.65e-20
C16185 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# V_LOW -2.78e-35
C16186 sky130_fd_sc_hd__dfbbn_1_46/Q_N V_GND -0.00252f
C16187 sky130_fd_sc_hd__conb_1_23/LO sky130_fd_sc_hd__inv_1_53/Y 0.0316f
C16188 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 1.63e-19
C16189 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# -0.00263f
C16190 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__dfbbn_1_7/a_941_21# -7.6e-19
C16191 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# -5.54e-21
C16192 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_47/Y 0.00419f
C16193 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 0.01f
C16194 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.66e-19
C16195 sky130_fd_sc_hd__dfbbn_1_32/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF3.Q 3.25e-19
C16196 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# sky130_fd_sc_hd__conb_1_35/HI 7.42e-20
C16197 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# Reset 3.01e-21
C16198 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_16_2/Y 0.535f
C16199 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 0.0232f
C16200 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0284f
C16201 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0232f
C16202 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0.00102f
C16203 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 2.57e-21
C16204 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# sky130_fd_sc_hd__inv_16_1/Y 1.93e-19
C16205 sky130_fd_sc_hd__conb_1_6/LO sky130_fd_sc_hd__conb_1_18/HI 1.42e-19
C16206 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# RISING_COUNTER.COUNT_SUB_DFF9.Q 4.17e-19
C16207 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.4e-20
C16208 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00604f
C16209 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0355f
C16210 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 8.1e-20
C16211 sky130_fd_sc_hd__fill_4_60/VPB V_GND 0.4f
C16212 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.0074f
C16213 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# FULL_COUNTER.COUNT_SUB_DFF16.Q 3.97e-20
C16214 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 2.75e-20
C16215 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_0/a_941_21# 1.9e-19
C16216 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# V_LOW 4.14e-20
C16217 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# FULL_COUNTER.COUNT_SUB_DFF5.Q 3.66e-19
C16218 sky130_fd_sc_hd__dfbbn_1_11/a_557_413# sky130_fd_sc_hd__inv_16_2/Y 5.67e-19
C16219 sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00149f
C16220 sky130_fd_sc_hd__dfbbn_1_8/a_1112_329# sky130_fd_sc_hd__inv_16_2/Y 0.001f
C16221 sky130_fd_sc_hd__dfbbn_1_25/a_581_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 4.53e-20
C16222 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# sky130_fd_sc_hd__conb_1_33/HI 0.00216f
C16223 sky130_fd_sc_hd__inv_16_2/Y FULL_COUNTER.COUNT_SUB_DFF18.Q 0.0294f
C16224 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# sky130_fd_sc_hd__conb_1_2/HI 0.00359f
C16225 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# -1.24e-20
C16226 sky130_fd_sc_hd__dfbbn_1_5/a_557_413# FULL_COUNTER.COUNT_SUB_DFF5.Q 0.00212f
C16227 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_39/A 4.48e-22
C16228 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# -0.00471f
C16229 sky130_fd_sc_hd__dfbbn_1_50/Q_N sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 1.18e-19
C16230 sky130_fd_sc_hd__conb_1_17/LO V_GND -6.11e-19
C16231 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 1.16e-19
C16232 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 2.87e-19
C16233 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 3.77e-19
C16234 sky130_fd_sc_hd__conb_1_48/HI sky130_fd_sc_hd__conb_1_36/HI 5e-20
C16235 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_93/A 0.112f
C16236 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__inv_1_100/Y 1.83e-19
C16237 sky130_fd_sc_hd__inv_1_107/Y V_GND 0.177f
C16238 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0147f
C16239 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0382f
C16240 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__inv_1_13/Y 0.0033f
C16241 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 1.52e-19
C16242 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# 5.77e-20
C16243 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 2.02e-20
C16244 sky130_fd_sc_hd__dfbbn_1_14/Q_N sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 7.72e-21
C16245 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# RISING_COUNTER.COUNT_SUB_DFF6.Q 8.29e-20
C16246 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__conb_1_45/HI 0.0172f
C16247 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 0.00249f
C16248 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0423f
C16249 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# V_LOW 0.00607f
C16250 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# V_LOW -0.308f
C16251 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 6.31e-21
C16252 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 3.23e-21
C16253 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# V_LOW 1.38e-19
C16254 sky130_fd_sc_hd__inv_1_107/Y sky130_fd_sc_hd__inv_1_106/Y 0.16f
C16255 sky130_fd_sc_hd__conb_1_44/HI sky130_fd_sc_hd__conb_1_45/HI 0.0291f
C16256 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# V_LOW 0.00607f
C16257 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_13/a_193_47# -0.0413f
C16258 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0326f
C16259 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# sky130_fd_sc_hd__inv_16_1/Y 0.0305f
C16260 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# V_LOW -6.44e-19
C16261 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__inv_16_0/Y 0.00303f
C16262 sky130_fd_sc_hd__dfbbn_1_49/Q_N FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.019f
C16263 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF11.Q 4.56e-21
C16264 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.00176f
C16265 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 4.43e-19
C16266 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0.00234f
C16267 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# sky130_fd_sc_hd__dfbbn_1_46/a_581_47# -7.91e-19
C16268 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.566f
C16269 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# V_LOW 0.00625f
C16270 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_119/Y 0.00317f
C16271 sky130_fd_sc_hd__conb_1_33/HI Reset 0.0894f
C16272 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 8.96e-20
C16273 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# V_GND -0.00501f
C16274 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# V_GND -0.0466f
C16275 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# sky130_fd_sc_hd__conb_1_22/HI 0.00113f
C16276 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__inv_1_62/Y 0.454f
C16277 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# V_LOW 0.0153f
C16278 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# sky130_fd_sc_hd__dfbbn_1_4/Q_N -4.33e-20
C16279 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__conb_1_28/LO 8.18e-19
C16280 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__dfbbn_1_2/a_473_413# -3.86e-20
C16281 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# sky130_fd_sc_hd__dfbbn_1_2/a_941_21# -1.03e-19
C16282 sky130_fd_sc_hd__dfbbn_1_49/Q_N V_LOW -0.00141f
C16283 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 0.0666f
C16284 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.131f
C16285 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 2.16f
C16286 sky130_fd_sc_hd__dfbbn_1_15/a_1112_329# V_GND 6.28e-19
C16287 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# V_GND 0.00529f
C16288 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# -9.32e-20
C16289 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 4.06e-21
C16290 sky130_fd_sc_hd__dfbbn_1_6/Q_N FULL_COUNTER.COUNT_SUB_DFF10.Q 2.07e-20
C16291 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_13/a_1672_329# 4.01e-19
C16292 sky130_fd_sc_hd__dfbbn_1_3/Q_N FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00128f
C16293 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# V_GND 7.9e-19
C16294 sky130_fd_sc_hd__dfbbn_1_31/a_1363_47# sky130_fd_sc_hd__conb_1_35/HI -2.65e-20
C16295 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_91/A 0.137f
C16296 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# sky130_fd_sc_hd__conb_1_45/HI 0.00274f
C16297 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# sky130_fd_sc_hd__dfbbn_1_39/Q_N 5.48e-20
C16298 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0.00135f
C16299 sky130_fd_sc_hd__conb_1_23/HI RISING_COUNTER.COUNT_SUB_DFF2.Q 1.08e-19
C16300 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__inv_1_10/Y 0.0139f
C16301 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.00881f
C16302 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.0549f
C16303 sky130_fd_sc_hd__conb_1_25/HI RISING_COUNTER.COUNT_SUB_DFF2.Q 0.402f
C16304 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0.00126f
C16305 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 2.65e-20
C16306 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 0.15f
C16307 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 1.52e-20
C16308 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# sky130_fd_sc_hd__conb_1_49/HI -5.09e-21
C16309 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# sky130_fd_sc_hd__inv_1_106/Y 2.67e-19
C16310 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# V_GND -0.00272f
C16311 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__inv_1_15/Y 3.81e-19
C16312 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_59/Y 0.251f
C16313 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# V_GND 0.00458f
C16314 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.325f
C16315 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.00307f
C16316 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0397f
C16317 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 2.23e-20
C16318 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF7.Q 9.47e-19
C16319 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# 4.54e-21
C16320 sky130_fd_sc_hd__dfbbn_1_17/Q_N V_LOW 1.99e-19
C16321 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# V_LOW 0.0059f
C16322 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# sky130_fd_sc_hd__inv_16_0/Y 1.74e-19
C16323 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# sky130_fd_sc_hd__inv_1_23/Y 1.88e-19
C16324 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 0.00332f
C16325 sky130_fd_sc_hd__inv_1_91/Y sky130_fd_sc_hd__inv_1_86/Y 0.108f
C16326 RISING_COUNTER.COUNT_SUB_DFF15.Q V_LOW 1.76f
C16327 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# sky130_fd_sc_hd__conb_1_33/HI 0.0047f
C16328 sky130_fd_sc_hd__dfbbn_1_39/a_1363_47# sky130_fd_sc_hd__conb_1_46/HI 4.08e-19
C16329 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 1.57e-20
C16330 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__dfbbn_1_37/a_581_47# -2.6e-20
C16331 sky130_fd_sc_hd__inv_1_9/Y FULL_COUNTER.COUNT_SUB_DFF2.Q 0.00399f
C16332 sky130_fd_sc_hd__conb_1_0/HI sky130_fd_sc_hd__inv_1_5/Y 6.8e-19
C16333 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__dfbbn_1_9/Q_N -4.97e-19
C16334 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 1.41e-19
C16335 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__inv_1_21/Y 3.98e-19
C16336 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 1.18e-20
C16337 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 9.56e-21
C16338 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__dfbbn_1_42/a_193_47# -0.11f
C16339 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# 1.75e-20
C16340 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# sky130_fd_sc_hd__inv_16_2/Y 0.0997f
C16341 sky130_fd_sc_hd__dfbbn_1_15/a_557_413# sky130_fd_sc_hd__inv_1_20/Y 8.17e-19
C16342 RISING_COUNTER.COUNT_SUB_DFF6.Q RISING_COUNTER.COUNT_SUB_DFF4.Q 3.29e-20
C16343 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF9.Q 6.62e-20
C16344 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_62/Y 0.135f
C16345 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_941_21# -0.00151f
C16346 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# -2.25e-19
C16347 sky130_fd_sc_hd__nand2_8_7/a_27_47# sky130_fd_sc_hd__inv_1_70/A 0.0288f
C16348 FULL_COUNTER.COUNT_SUB_DFF15.Q FULL_COUNTER.COUNT_SUB_DFF0.Q 0.104f
C16349 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# V_GND 0.00337f
C16350 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# sky130_fd_sc_hd__inv_1_11/Y 0.00196f
C16351 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_105/Y 0.0531f
C16352 sky130_fd_sc_hd__dfbbn_1_6/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 2.44e-20
C16353 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0147f
C16354 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 7.88e-19
C16355 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# sky130_fd_sc_hd__inv_1_99/Y 2.87e-20
C16356 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# FULL_COUNTER.COUNT_SUB_DFF11.Q 4.36e-20
C16357 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# sky130_fd_sc_hd__conb_1_45/HI 0.00526f
C16358 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.0514f
C16359 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# sky130_fd_sc_hd__inv_1_17/Y 2.22e-19
C16360 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 6.96e-20
C16361 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# sky130_fd_sc_hd__conb_1_8/HI 1.36e-19
C16362 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.11e-19
C16363 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 6.12e-19
C16364 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 4.61e-21
C16365 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 3.71e-20
C16366 sky130_fd_sc_hd__dfbbn_1_13/a_1159_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00178f
C16367 sky130_fd_sc_hd__conb_1_47/HI FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.0064f
C16368 RISING_COUNTER.COUNT_SUB_DFF11.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0632f
C16369 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__inv_16_0/Y 0.00327f
C16370 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# V_LOW -0.315f
C16371 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 7.06e-19
C16372 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__conb_1_50/LO 0.0144f
C16373 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_108/Y 8.09e-19
C16374 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00223f
C16375 sky130_fd_sc_hd__conb_1_20/HI V_GND 0.21f
C16376 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF4.Q 0.402f
C16377 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 1.21e-19
C16378 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 1.21e-19
C16379 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 1.81e-19
C16380 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 1.81e-19
C16381 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# sky130_fd_sc_hd__inv_1_17/Y 0.00225f
C16382 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# V_GND -0.00493f
C16383 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# V_GND 1.82e-19
C16384 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# sky130_fd_sc_hd__conb_1_22/HI 1.39e-19
C16385 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_12/HI 6.44e-19
C16386 sky130_fd_sc_hd__dfbbn_1_44/a_1340_413# V_LOW 2.94e-20
C16387 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# sky130_fd_sc_hd__inv_1_105/Y 0.00458f
C16388 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__dfbbn_1_2/a_1340_413# -2.57e-20
C16389 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_16_1/Y 2.72e-19
C16390 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# 0.00195f
C16391 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.157f
C16392 sky130_fd_sc_hd__dfbbn_1_4/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 5.64e-19
C16393 sky130_fd_sc_hd__dfbbn_1_31/a_1672_329# V_GND 2.56e-19
C16394 sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF9.Q 0.00434f
C16395 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# sky130_fd_sc_hd__dfbbn_1_7/Q_N -4.33e-20
C16396 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# FALLING_COUNTER.COUNT_SUB_DFF1.Q 1.04e-20
C16397 RISING_COUNTER.COUNT_SUB_DFF9.Q sky130_fd_sc_hd__conb_1_28/HI 2.51e-19
C16398 sky130_fd_sc_hd__conb_1_31/HI sky130_fd_sc_hd__inv_1_60/Y 1.82e-20
C16399 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# V_GND 3.08e-19
C16400 sky130_fd_sc_hd__conb_1_6/HI V_LOW 0.168f
C16401 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# V_LOW 2.25e-19
C16402 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 0.0011f
C16403 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# V_GND 0.00646f
C16404 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# sky130_fd_sc_hd__dfbbn_1_38/a_381_47# -3.79e-20
C16405 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_1112_329# -4.66e-20
C16406 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# CLOCK_GEN.SR_Op.Q 1.86e-19
C16407 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# sky130_fd_sc_hd__conb_1_46/HI 9.05e-20
C16408 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_48/a_1340_413# 1.02e-19
C16409 sky130_fd_sc_hd__conb_1_8/LO sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 9.17e-19
C16410 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 5.49e-20
C16411 sky130_fd_sc_hd__nand3_1_2/Y sky130_fd_sc_hd__inv_16_1/Y 1.15e-20
C16412 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.29e-19
C16413 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 1.04e-20
C16414 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 8.03e-21
C16415 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# sky130_fd_sc_hd__dfbbn_1_50/a_1112_329# -4.66e-20
C16416 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# sky130_fd_sc_hd__dfbbn_1_50/a_381_47# -3.79e-20
C16417 sky130_fd_sc_hd__dfbbn_1_38/a_1159_47# sky130_fd_sc_hd__conb_1_49/HI 2.06e-20
C16418 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF15.Q 7.11e-20
C16419 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# V_GND -0.00304f
C16420 FALLING_COUNTER.COUNT_SUB_DFF4.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.0295f
C16421 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# sky130_fd_sc_hd__inv_1_59/Y 0.00388f
C16422 sky130_fd_sc_hd__dfbbn_1_44/a_1159_47# V_GND 8.02e-19
C16423 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 1.22e-19
C16424 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.00399f
C16425 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 1.07e-19
C16426 sky130_fd_sc_hd__dfbbn_1_34/Q_N FALLING_COUNTER.COUNT_SUB_DFF11.Q 0.0215f
C16427 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# sky130_fd_sc_hd__conb_1_42/HI 2.78e-19
C16428 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 0.00923f
C16429 sky130_fd_sc_hd__dfbbn_1_19/a_891_329# FULL_COUNTER.COUNT_SUB_DFF2.Q 1.08e-19
C16430 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF2.Q 3.66e-20
C16431 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.00528f
C16432 sky130_fd_sc_hd__dfbbn_1_19/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00835f
C16433 sky130_fd_sc_hd__conb_1_40/LO V_GND -0.00266f
C16434 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# RISING_COUNTER.COUNT_SUB_DFF4.Q 0.0297f
C16435 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 5.1e-19
C16436 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_941_21# -0.00248f
C16437 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# -7.77e-19
C16438 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 3.41e-19
C16439 sky130_fd_sc_hd__dfbbn_1_51/a_1112_329# V_GND 7.66e-19
C16440 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_381_47# -0.00441f
C16441 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# sky130_fd_sc_hd__inv_1_23/Y 4.42e-19
C16442 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_94/A 1.31e-19
C16443 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# sky130_fd_sc_hd__inv_16_2/Y 4.71e-20
C16444 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 5.94e-19
C16445 FULL_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__conb_1_5/HI 0.0131f
C16446 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 8.14e-19
C16447 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# sky130_fd_sc_hd__inv_1_10/Y 4.23e-21
C16448 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF9.Q 1.81e-20
C16449 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00814f
C16450 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0.00246f
C16451 sky130_fd_sc_hd__dfbbn_1_7/a_1672_329# sky130_fd_sc_hd__inv_16_2/Y 2.4e-20
C16452 FULL_COUNTER.COUNT_SUB_DFF10.Q V_GND 3.52f
C16453 sky130_fd_sc_hd__conb_1_22/HI sky130_fd_sc_hd__inv_1_53/Y 0.566f
C16454 sky130_fd_sc_hd__conb_1_49/HI sky130_fd_sc_hd__inv_16_1/Y 0.201f
C16455 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 2.29e-19
C16456 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# sky130_fd_sc_hd__inv_1_63/Y 9.37e-19
C16457 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF9.Q 1.72e-20
C16458 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# sky130_fd_sc_hd__dfbbn_1_3/a_473_413# -3.06e-20
C16459 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# sky130_fd_sc_hd__dfbbn_1_3/a_647_21# -6.43e-20
C16460 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# -1.63e-19
C16461 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# sky130_fd_sc_hd__dfbbn_1_23/a_1672_329# -7.17e-20
C16462 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__inv_1_54/Y 4.23e-21
C16463 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# sky130_fd_sc_hd__inv_1_60/Y 4.94e-20
C16464 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# RISING_COUNTER.COUNT_SUB_DFF4.Q 2.22e-19
C16465 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# V_GND 0.00179f
C16466 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_2_0/Y 2.54e-20
C16467 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# sky130_fd_sc_hd__inv_1_11/Y 7.95e-19
C16468 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 1.76e-20
C16469 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0475f
C16470 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 7.52e-22
C16471 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# -7.77e-19
C16472 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_941_21# -0.00153f
C16473 sky130_fd_sc_hd__inv_1_104/Y FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.401f
C16474 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.0215f
C16475 sky130_fd_sc_hd__inv_16_0/Y sky130_fd_sc_hd__conb_1_28/HI 0.484f
C16476 sky130_fd_sc_hd__conb_1_10/HI sky130_fd_sc_hd__conb_1_18/HI 3.25e-19
C16477 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# V_LOW 0.0169f
C16478 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# -2.37e-19
C16479 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__dfbbn_1_47/a_941_21# -0.00139f
C16480 FULL_COUNTER.COUNT_SUB_DFF17.Q V_LOW 0.463f
C16481 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0167f
C16482 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00101f
C16483 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 1.1e-20
C16484 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00319f
C16485 sky130_fd_sc_hd__conb_1_50/LO RISING_COUNTER.COUNT_SUB_DFF7.Q 3.89e-20
C16486 sky130_fd_sc_hd__inv_1_64/Y sky130_fd_sc_hd__inv_1_94/Y 0.0398f
C16487 sky130_fd_sc_hd__conb_1_51/HI V_GND 0.0926f
C16488 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 7.21e-20
C16489 sky130_fd_sc_hd__conb_1_41/LO sky130_fd_sc_hd__conb_1_40/HI 1.82e-20
C16490 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__inv_16_0/Y 0.026f
C16491 sky130_fd_sc_hd__inv_1_89/Y sky130_fd_sc_hd__inv_1_83/Y 0.364f
C16492 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 4.43e-20
C16493 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 3.24e-19
C16494 sky130_fd_sc_hd__inv_1_71/Y sky130_fd_sc_hd__inv_1_70/Y 0.00381f
C16495 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# sky130_fd_sc_hd__inv_1_5/Y 0.00645f
C16496 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF12.Q 3.27e-21
C16497 sky130_fd_sc_hd__conb_1_11/LO FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00281f
C16498 sky130_fd_sc_hd__dfbbn_1_51/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF0.Q 4.6e-20
C16499 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 1.08e-19
C16500 sky130_fd_sc_hd__dfbbn_1_31/a_1340_413# FALLING_COUNTER.COUNT_SUB_DFF4.Q 2.59e-19
C16501 FULL_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_12/Y 0.00696f
C16502 sky130_fd_sc_hd__inv_1_11/Y FULL_COUNTER.COUNT_SUB_DFF11.Q 0.14f
C16503 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# sky130_fd_sc_hd__inv_1_90/Y 0.00488f
C16504 sky130_fd_sc_hd__inv_1_80/A sky130_fd_sc_hd__inv_1_68/A 9.24e-20
C16505 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# sky130_fd_sc_hd__conb_1_25/HI 4.95e-19
C16506 sky130_fd_sc_hd__dfbbn_1_11/a_891_329# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00138f
C16507 sky130_fd_sc_hd__conb_1_38/HI sky130_fd_sc_hd__inv_1_76/A 3.23e-20
C16508 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_9/Y 0.107f
C16509 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# FULL_COUNTER.COUNT_SUB_DFF5.Q 2.38e-20
C16510 sky130_fd_sc_hd__dfbbn_1_22/Q_N V_GND 0.00216f
C16511 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.98e-20
C16512 sky130_fd_sc_hd__dfbbn_1_30/a_557_413# V_GND 2.09e-19
C16513 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__inv_16_2/Y 0.0419f
C16514 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# V_LOW 0.00616f
C16515 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# sky130_fd_sc_hd__dfbbn_1_17/a_381_47# -0.00171f
C16516 sky130_fd_sc_hd__dfbbn_1_45/Q_N V_GND -0.00803f
C16517 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 1.14e-19
C16518 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_15/a_1159_47# 3.16e-19
C16519 sky130_fd_sc_hd__dfbbn_1_19/a_1672_329# V_GND 2.85e-19
C16520 sky130_fd_sc_hd__conb_1_14/HI sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 7.9e-20
C16521 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__inv_16_0/Y 0.00162f
C16522 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# sky130_fd_sc_hd__inv_16_1/Y 1.29e-19
C16523 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 9.73e-21
C16524 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 3.68e-21
C16525 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 5.11e-21
C16526 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 9.23e-20
C16527 sky130_fd_sc_hd__dfbbn_1_2/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.66e-19
C16528 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# sky130_fd_sc_hd__dfbbn_1_0/a_557_413# -0.0012f
C16529 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# -0.00736f
C16530 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 0.00516f
C16531 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_1/a_473_413# 6.67e-20
C16532 sky130_fd_sc_hd__dfbbn_1_45/Q_N sky130_fd_sc_hd__inv_1_106/Y 0.00355f
C16533 sky130_fd_sc_hd__dfbbn_1_18/Q_N V_GND -0.00769f
C16534 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__inv_1_19/Y 0.00551f
C16535 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# 8.24e-19
C16536 sky130_fd_sc_hd__dfbbn_1_9/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.0254f
C16537 sky130_fd_sc_hd__dfbbn_1_46/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.57e-19
C16538 sky130_fd_sc_hd__dfbbn_1_3/a_557_413# sky130_fd_sc_hd__inv_16_2/Y 4.66e-21
C16539 sky130_fd_sc_hd__dfbbn_1_40/Q_N FALLING_COUNTER.COUNT_SUB_DFF7.Q 5.4e-21
C16540 sky130_fd_sc_hd__dfbbn_1_35/a_557_413# V_GND 5.55e-19
C16541 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 1.11e-19
C16542 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# -1.66e-19
C16543 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_40/A 0.00914f
C16544 sky130_fd_sc_hd__dfbbn_1_7/Q_N sky130_fd_sc_hd__inv_1_23/Y 0.0203f
C16545 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__conb_1_40/HI 0.00189f
C16546 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1672_329# -1.44e-20
C16547 FULL_COUNTER.COUNT_SUB_DFF19.Q V_GND 2.73f
C16548 sky130_fd_sc_hd__nand2_8_9/a_27_47# sky130_fd_sc_hd__inv_1_70/Y 1.02e-19
C16549 sky130_fd_sc_hd__inv_1_81/Y sky130_fd_sc_hd__inv_1_92/Y 8.79e-20
C16550 RISING_COUNTER.COUNT_SUB_DFF14.Q RISING_COUNTER.COUNT_SUB_DFF13.Q 0.166f
C16551 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 5.77e-22
C16552 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF11.Q 0.00758f
C16553 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 4.8e-19
C16554 sky130_fd_sc_hd__nand3_1_0/Y sky130_fd_sc_hd__inv_1_72/A 0.00112f
C16555 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_75/Y 0.00422f
C16556 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# -3.48e-20
C16557 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# sky130_fd_sc_hd__dfbbn_1_43/a_891_329# -2.2e-20
C16558 sky130_fd_sc_hd__conb_1_8/HI sky130_fd_sc_hd__dfbbn_1_5/a_1159_47# -0.00236f
C16559 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# CLOCK_GEN.SR_Op.Q 3.49e-19
C16560 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF3.Q 1.37f
C16561 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__conb_1_12/LO 1.64e-21
C16562 sky130_fd_sc_hd__conb_1_37/LO V_GND 0.00248f
C16563 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 1.8e-20
C16564 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_34/a_1112_329# 0.00408f
C16565 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 5.99e-20
C16566 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 3.06e-21
C16567 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# sky130_fd_sc_hd__conb_1_4/LO 1.53e-19
C16568 sky130_fd_sc_hd__conb_1_39/HI sky130_fd_sc_hd__conb_1_41/HI 0.00375f
C16569 sky130_fd_sc_hd__inv_1_111/Y RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0915f
C16570 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 6.89e-19
C16571 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 8.98e-19
C16572 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 3.03e-21
C16573 sky130_fd_sc_hd__inv_1_21/Y FULL_COUNTER.COUNT_SUB_DFF13.Q 4.64e-19
C16574 sky130_fd_sc_hd__dfbbn_1_25/Q_N V_GND -9.87e-19
C16575 sky130_fd_sc_hd__dfbbn_1_4/Q_N sky130_fd_sc_hd__inv_1_11/Y 5.04e-21
C16576 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1_0/Y 0.00286f
C16577 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# -7.17e-20
C16578 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_27/a_791_47# -2.22e-34
C16579 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# -1.66e-19
C16580 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 5.74e-19
C16581 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00245f
C16582 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# V_LOW 5.11e-19
C16583 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__conb_1_17/HI 0.0485f
C16584 sky130_fd_sc_hd__conb_1_48/LO V_GND -0.00351f
C16585 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# FULL_COUNTER.COUNT_SUB_DFF11.Q 2.73e-19
C16586 FALLING_COUNTER.COUNT_SUB_DFF2.Q sky130_fd_sc_hd__dfbbn_1_32/a_557_413# 2.83e-19
C16587 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# V_LOW 0.00836f
C16588 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# -1.66e-19
C16589 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0102f
C16590 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# sky130_fd_sc_hd__conb_1_8/HI 6.67e-20
C16591 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# sky130_fd_sc_hd__conb_1_6/HI 0.0336f
C16592 sky130_fd_sc_hd__conb_1_21/LO V_GND -0.006f
C16593 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 0.0102f
C16594 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 0.00127f
C16595 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 8.32e-19
C16596 sky130_fd_sc_hd__nand2_1_5/Y sky130_fd_sc_hd__inv_1_76/A 2.35e-20
C16597 sky130_fd_sc_hd__conb_1_48/LO sky130_fd_sc_hd__inv_1_106/Y 0.0412f
C16598 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__inv_1_99/Y 1.24e-21
C16599 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.54e-19
C16600 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0.105f
C16601 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 4.15e-19
C16602 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# RISING_COUNTER.COUNT_SUB_DFF2.Q 8.41e-21
C16603 sky130_fd_sc_hd__dfbbn_1_21/a_1363_47# sky130_fd_sc_hd__conb_1_25/HI 4.16e-19
C16604 sky130_fd_sc_hd__conb_1_44/LO sky130_fd_sc_hd__conb_1_49/LO 0.236f
C16605 FULL_COUNTER.COUNT_SUB_DFF5.Q sky130_fd_sc_hd__conb_1_5/HI 9.51e-20
C16606 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# V_GND 0.0043f
C16607 RISING_COUNTER.COUNT_SUB_DFF9.Q V_GND 0.924f
C16608 sky130_fd_sc_hd__inv_1_108/Y sky130_fd_sc_hd__inv_1_59/Y 2.37e-20
C16609 FULL_COUNTER.COUNT_SUB_DFF13.Q FULL_COUNTER.COUNT_SUB_DFF18.Q 6.81e-20
C16610 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 4.35e-22
C16611 sky130_fd_sc_hd__conb_1_30/LO sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 1.87e-22
C16612 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00829f
C16613 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# sky130_fd_sc_hd__inv_16_2/Y 0.00478f
C16614 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF3.Q 0.0206f
C16615 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# V_LOW 8.06e-19
C16616 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.76e-20
C16617 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_17/a_1672_329# -1.44e-20
C16618 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__conb_1_31/HI 3.14e-20
C16619 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00426f
C16620 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# 0.00104f
C16621 sky130_fd_sc_hd__dfbbn_1_40/a_1112_329# FALLING_COUNTER.COUNT_SUB_DFF8.Q 1.97e-19
C16622 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# sky130_fd_sc_hd__conb_1_24/HI 2.46e-20
C16623 FULL_COUNTER.COUNT_SUB_DFF19.Q sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 2.1e-20
C16624 sky130_fd_sc_hd__nand2_8_2/a_27_47# sky130_fd_sc_hd__nand2_1_2/A 5.43e-19
C16625 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# V_GND 0.035f
C16626 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# -5.42e-19
C16627 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.29e-19
C16628 sky130_fd_sc_hd__inv_1_31/A V_SENSE 0.0487f
C16629 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_108/Y 4.81e-21
C16630 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# sky130_fd_sc_hd__inv_1_19/Y 1.44e-21
C16631 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_37/Q_N 0.0024f
C16632 sky130_fd_sc_hd__conb_1_14/HI FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00186f
C16633 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0359f
C16634 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__inv_16_2/Y 0.0738f
C16635 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# sky130_fd_sc_hd__conb_1_5/HI 7.79e-19
C16636 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__conb_1_27/HI 3.41e-19
C16637 sky130_fd_sc_hd__conb_1_20/HI RISING_COUNTER.COUNT_SUB_DFF12.Q 0.0257f
C16638 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 5.59e-20
C16639 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# sky130_fd_sc_hd__conb_1_28/HI 9.75e-20
C16640 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# sky130_fd_sc_hd__inv_16_2/Y 0.0172f
C16641 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 0.00116f
C16642 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# sky130_fd_sc_hd__inv_1_50/A 2e-19
C16643 sky130_fd_sc_hd__conb_1_25/HI sky130_fd_sc_hd__conb_1_26/LO 0.0849f
C16644 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# -3.46e-20
C16645 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__nand2_8_3/a_27_47# 1.26e-21
C16646 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF7.Q 2.81e-20
C16647 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_12/a_581_47# 4.29e-20
C16648 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 7.04e-19
C16649 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 7.01e-19
C16650 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 4.62e-20
C16651 sky130_fd_sc_hd__inv_16_0/Y V_GND 4.09f
C16652 sky130_fd_sc_hd__dfbbn_1_43/Q_N sky130_fd_sc_hd__inv_1_60/Y 1.7e-19
C16653 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__inv_1_56/Y 1.62e-19
C16654 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# sky130_fd_sc_hd__conb_1_23/HI -0.00234f
C16655 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# sky130_fd_sc_hd__inv_16_2/Y 0.0191f
C16656 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 1.51e-20
C16657 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 1.09e-19
C16658 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 1.14e-20
C16659 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 3.21e-20
C16660 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 1.25e-20
C16661 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__conb_1_19/LO 3.46e-20
C16662 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0.00491f
C16663 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.18e-21
C16664 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# sky130_fd_sc_hd__conb_1_25/HI 0.0181f
C16665 sky130_fd_sc_hd__dfbbn_1_12/Q_N FULL_COUNTER.COUNT_SUB_DFF16.Q 0.0274f
C16666 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00478f
C16667 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__inv_1_90/Y 0.053f
C16668 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# RISING_COUNTER.COUNT_SUB_DFF1.Q 1.33e-22
C16669 Reset sky130_fd_sc_hd__inv_1_99/Y 2.85e-20
C16670 sky130_fd_sc_hd__inv_1_109/Y FALLING_COUNTER.COUNT_SUB_DFF9.Q 8.95e-19
C16671 RISING_COUNTER.COUNT_SUB_DFF7.Q RISING_COUNTER.COUNT_SUB_DFF6.Q 0.244f
C16672 sky130_fd_sc_hd__inv_1_62/Y RISING_COUNTER.COUNT_SUB_DFF5.Q 5.49e-20
C16673 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.51e-19
C16674 FULL_COUNTER.COUNT_SUB_DFF17.Q sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 0.0511f
C16675 sky130_fd_sc_hd__dfbbn_1_14/a_557_413# FULL_COUNTER.COUNT_SUB_DFF8.Q 4.43e-19
C16676 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# sky130_fd_sc_hd__inv_1_101/Y 0.0037f
C16677 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 1.8e-20
C16678 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0115f
C16679 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_38/LO 6.52e-20
C16680 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 2.55e-19
C16681 FULL_COUNTER.COUNT_SUB_DFF15.Q RISING_COUNTER.COUNT_SUB_DFF0.Q 0.00132f
C16682 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF4.Q 3.95e-20
C16683 sky130_fd_sc_hd__conb_1_16/HI sky130_fd_sc_hd__inv_1_22/Y 2.93e-20
C16684 sky130_fd_sc_hd__nand3_1_2/Y FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00219f
C16685 sky130_fd_sc_hd__dfbbn_1_47/a_891_329# CLOCK_GEN.SR_Op.Q 0.00283f
C16686 sky130_fd_sc_hd__dfbbn_1_21/a_891_329# V_LOW -0.00121f
C16687 sky130_fd_sc_hd__inv_1_89/Y V_LOW 0.0462f
C16688 sky130_fd_sc_hd__inv_1_83/Y sky130_fd_sc_hd__inv_1_95/A 9.39e-19
C16689 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF9.Q 0.0037f
C16690 sky130_fd_sc_hd__dfbbn_1_4/a_891_329# FULL_COUNTER.COUNT_SUB_DFF10.Q 8.56e-19
C16691 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# V_GND 0.00281f
C16692 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# sky130_fd_sc_hd__inv_1_54/Y 0.00352f
C16693 sky130_fd_sc_hd__dfbbn_1_16/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 6.69e-20
C16694 sky130_fd_sc_hd__inv_1_91/Y V_GND 0.117f
C16695 sky130_fd_sc_hd__inv_1_19/Y sky130_fd_sc_hd__inv_16_2/Y 0.0156f
C16696 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 3.76e-19
C16697 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# FULL_COUNTER.COUNT_SUB_DFF13.Q 4.46e-20
C16698 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0.0113f
C16699 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 8.77e-20
C16700 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.00174f
C16701 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 5.27e-20
C16702 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 3.21e-19
C16703 FULL_COUNTER.COUNT_SUB_DFF14.Q FULL_COUNTER.COUNT_SUB_DFF5.Q 4.16e-20
C16704 sky130_fd_sc_hd__nand3_1_2/Y V_LOW 0.519f
C16705 sky130_fd_sc_hd__dfbbn_1_21/a_1112_329# sky130_fd_sc_hd__conb_1_26/HI 0.00107f
C16706 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 3.24e-20
C16707 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# sky130_fd_sc_hd__inv_16_0/Y 1.42e-19
C16708 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF16.Q 0.00503f
C16709 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__inv_1_18/Y 2.32e-20
C16710 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# sky130_fd_sc_hd__inv_16_1/Y 0.0385f
C16711 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# V_GND 0.00366f
C16712 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# sky130_fd_sc_hd__conb_1_6/HI 0.00217f
C16713 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0313f
C16714 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 0.0167f
C16715 sky130_fd_sc_hd__conb_1_3/HI sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.0134f
C16716 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__conb_1_46/HI 2.04e-20
C16717 RISING_COUNTER.COUNT_SUB_DFF8.Q sky130_fd_sc_hd__dfbbn_1_24/Q_N 0.00266f
C16718 sky130_fd_sc_hd__dfbbn_1_51/Q_N FALLING_COUNTER.COUNT_SUB_DFF4.Q 4.33e-20
C16719 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# CLOCK_GEN.SR_Op.Q 1.96e-20
C16720 sky130_fd_sc_hd__inv_1_39/Y V_GND 0.137f
C16721 sky130_fd_sc_hd__conb_1_1/HI FULL_COUNTER.COUNT_SUB_DFF4.Q 2.51e-19
C16722 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# sky130_fd_sc_hd__conb_1_22/HI 6.28e-20
C16723 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0409f
C16724 sky130_fd_sc_hd__conb_1_44/HI FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0915f
C16725 sky130_fd_sc_hd__conb_1_50/HI sky130_fd_sc_hd__dfbbn_1_43/a_557_413# 5.03e-19
C16726 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# V_GND 0.00835f
C16727 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 0.0039f
C16728 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_93/Y 0.00406f
C16729 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF7.Q 0.0102f
C16730 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# sky130_fd_sc_hd__inv_16_0/Y 0.0349f
C16731 sky130_fd_sc_hd__conb_1_7/LO sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 3.6e-21
C16732 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# sky130_fd_sc_hd__inv_1_99/Y 0.00992f
C16733 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 3.48e-19
C16734 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_71/A 0.0022f
C16735 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 2.56e-21
C16736 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# sky130_fd_sc_hd__conb_1_28/HI 2.6e-19
C16737 sky130_fd_sc_hd__conb_1_18/LO sky130_fd_sc_hd__conb_1_18/HI 0.0132f
C16738 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 4.41e-19
C16739 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# sky130_fd_sc_hd__inv_16_2/Y 0.0129f
C16740 sky130_fd_sc_hd__conb_1_49/HI V_LOW 0.125f
C16741 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 8.48e-19
C16742 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0.00116f
C16743 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0.00124f
C16744 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__dfbbn_1_50/a_647_21# 1.62e-19
C16745 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_941_21# -0.0128f
C16746 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# -2.3e-19
C16747 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# -0.00124f
C16748 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# sky130_fd_sc_hd__dfbbn_1_41/a_557_413# -3.67e-20
C16749 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_6/Y 0.0658f
C16750 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# sky130_fd_sc_hd__inv_16_2/Y 0.00343f
C16751 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# FULL_COUNTER.COUNT_SUB_DFF4.Q 7.71e-21
C16752 RISING_COUNTER.COUNT_SUB_DFF10.Q sky130_fd_sc_hd__conb_1_30/HI 0.449f
C16753 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0265f
C16754 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_18/HI 9.55e-20
C16755 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# sky130_fd_sc_hd__inv_1_98/Y 0.00224f
C16756 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# V_GND 0.00685f
C16757 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF3.Q 2.55e-22
C16758 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# sky130_fd_sc_hd__nand2_1_0/Y 6.56e-21
C16759 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# sky130_fd_sc_hd__conb_1_18/HI -1.14e-20
C16760 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# V_GND 0.0196f
C16761 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__conb_1_17/HI 3.34e-21
C16762 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_37/HI 0.0112f
C16763 FULL_COUNTER.COUNT_SUB_DFF4.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 7.64e-20
C16764 sky130_fd_sc_hd__dfbbn_1_27/a_1159_47# sky130_fd_sc_hd__conb_1_23/HI -0.00265f
C16765 sky130_fd_sc_hd__dfbbn_1_18/a_581_47# sky130_fd_sc_hd__inv_16_2/Y 0.00167f
C16766 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# V_GND 0.0148f
C16767 sky130_fd_sc_hd__conb_1_43/HI sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 1.38e-20
C16768 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 0.028f
C16769 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_27/a_1672_329# 3.31e-19
C16770 sky130_fd_sc_hd__inv_1_93/Y V_GND 0.00809f
C16771 sky130_fd_sc_hd__dfbbn_1_47/a_1159_47# sky130_fd_sc_hd__conb_1_25/HI -0.00259f
C16772 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_105/Y 0.425f
C16773 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_106/Y -0.00323f
C16774 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_647_21# -0.00123f
C16775 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_16/HI 8.2e-21
C16776 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_12/a_557_413# 0.00149f
C16777 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# sky130_fd_sc_hd__conb_1_12/HI 5.85e-19
C16778 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF13.Q 0.0307f
C16779 FULL_COUNTER.COUNT_SUB_DFF19.Q RISING_COUNTER.COUNT_SUB_DFF12.Q 4.39e-21
C16780 FULL_COUNTER.COUNT_SUB_DFF7.Q FULL_COUNTER.COUNT_SUB_DFF11.Q 5.93e-20
C16781 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# sky130_fd_sc_hd__dfbbn_1_15/a_891_329# -2.2e-20
C16782 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# -9.65e-20
C16783 FALLING_COUNTER.COUNT_SUB_DFF3.Q FALLING_COUNTER.COUNT_SUB_DFF5.Q 6.05e-19
C16784 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__conb_1_41/LO 8.81e-20
C16785 sky130_fd_sc_hd__inv_1_94/Y Reset 0.0093f
C16786 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_1/a_473_413# 0.0211f
C16787 sky130_fd_sc_hd__conb_1_2/HI sky130_fd_sc_hd__conb_1_5/HI 1.28e-22
C16788 sky130_fd_sc_hd__conb_1_41/HI V_GND 0.226f
C16789 FULL_COUNTER.COUNT_SUB_DFF12.Q V_LOW 0.623f
C16790 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 5.8e-21
C16791 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 5.66e-19
C16792 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# sky130_fd_sc_hd__conb_1_22/HI -1.32e-19
C16793 FULL_COUNTER.COUNT_SUB_DFF3.Q FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0922f
C16794 sky130_fd_sc_hd__dfbbn_1_39/Q_N V_GND -0.00219f
C16795 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_647_21# -0.00392f
C16796 RISING_COUNTER.COUNT_SUB_DFF11.Q V_LOW 1.75f
C16797 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF14.Q 4.65e-21
C16798 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF6.Q 1.69e-20
C16799 sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# sky130_fd_sc_hd__inv_1_54/Y 1.07e-21
C16800 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# sky130_fd_sc_hd__conb_1_16/HI 7.79e-19
C16801 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__inv_1_59/Y 0.303f
C16802 sky130_fd_sc_hd__conb_1_35/HI sky130_fd_sc_hd__inv_16_1/Y 0.0583f
C16803 sky130_fd_sc_hd__dfbbn_1_37/a_891_329# V_LOW 2.26e-20
C16804 sky130_fd_sc_hd__dfbbn_1_25/Q_N RISING_COUNTER.COUNT_SUB_DFF12.Q 0.00185f
C16805 sky130_fd_sc_hd__dfbbn_1_10/a_557_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.23e-19
C16806 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# V_LOW 0.00538f
C16807 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__dfbbn_1_20/a_473_413# 0.00656f
C16808 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# sky130_fd_sc_hd__conb_1_12/HI -4.02e-19
C16809 sky130_fd_sc_hd__dfbbn_1_48/a_1159_47# sky130_fd_sc_hd__inv_16_0/Y 4.12e-19
C16810 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 9.27e-19
C16811 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 7.88e-21
C16812 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 7.71e-22
C16813 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# V_LOW -0.00237f
C16814 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# sky130_fd_sc_hd__inv_1_102/Y 3.62e-19
C16815 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# -6.29e-19
C16816 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# sky130_fd_sc_hd__dfbbn_1_24/a_557_413# -3.67e-20
C16817 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# sky130_fd_sc_hd__dfbbn_1_24/a_891_329# -2.46e-19
C16818 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.00336f
C16819 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# sky130_fd_sc_hd__inv_16_1/Y 0.054f
C16820 sky130_fd_sc_hd__inv_1_104/Y sky130_fd_sc_hd__inv_1_110/Y 3.24e-19
C16821 sky130_fd_sc_hd__inv_1_64/A sky130_fd_sc_hd__inv_1_86/Y 7.23e-20
C16822 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__inv_1_103/Y 0.0499f
C16823 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF0.Q 0.00134f
C16824 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 1.65e-19
C16825 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 4.56e-21
C16826 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# FALLING_COUNTER.COUNT_SUB_DFF5.Q 2.97e-22
C16827 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_4/a_1340_413# 2.75e-19
C16828 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF14.Q 4.56e-20
C16829 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# RISING_COUNTER.COUNT_SUB_DFF6.Q 3.6e-20
C16830 sky130_fd_sc_hd__dfbbn_1_47/Q_N RISING_COUNTER.COUNT_SUB_DFF0.Q 0.0364f
C16831 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# FULL_COUNTER.COUNT_SUB_DFF8.Q 2.07e-21
C16832 sky130_fd_sc_hd__conb_1_29/HI sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 0.00867f
C16833 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_647_21# -0.00157f
C16834 sky130_fd_sc_hd__dfbbn_1_2/a_1112_329# V_LOW 4.8e-20
C16835 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_57/Y 1.79e-19
C16836 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# V_GND 0.00186f
C16837 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.0378f
C16838 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.82e-19
C16839 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# sky130_fd_sc_hd__inv_1_99/Y 0.0054f
C16840 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.15f
C16841 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# V_GND 0.00418f
C16842 sky130_fd_sc_hd__dfbbn_1_38/a_557_413# V_LOW 3.56e-20
C16843 sky130_fd_sc_hd__dfbbn_1_45/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF7.Q 1.05e-20
C16844 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# sky130_fd_sc_hd__inv_16_0/Y 0.0351f
C16845 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# FULL_COUNTER.COUNT_SUB_DFF2.Q 0.1f
C16846 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00857f
C16847 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# sky130_fd_sc_hd__inv_1_99/Y 0.0306f
C16848 sky130_fd_sc_hd__dfbbn_1_50/a_557_413# V_LOW 3.56e-20
C16849 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__conb_1_35/HI 0.0243f
C16850 sky130_fd_sc_hd__dfbbn_1_23/a_557_413# V_GND 1.48e-19
C16851 sky130_fd_sc_hd__dfbbn_1_42/Q_N sky130_fd_sc_hd__conb_1_28/HI 5.05e-19
C16852 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 1.06e-20
C16853 sky130_fd_sc_hd__dfbbn_1_15/Q_N sky130_fd_sc_hd__inv_16_2/Y 0.00558f
C16854 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 3.95e-19
C16855 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0.0105f
C16856 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 4.7e-20
C16857 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 7.23e-19
C16858 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 4.74e-20
C16859 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 2.44e-20
C16860 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# sky130_fd_sc_hd__conb_1_40/HI 0.00508f
C16861 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 7.9e-19
C16862 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# sky130_fd_sc_hd__conb_1_9/HI 1.52e-22
C16863 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# RISING_COUNTER.COUNT_SUB_DFF10.Q 1.24e-20
C16864 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0235f
C16865 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# sky130_fd_sc_hd__dfbbn_1_33/a_1672_329# -5.16e-20
C16866 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# -1.66e-19
C16867 sky130_fd_sc_hd__inv_1_46/A sky130_fd_sc_hd__inv_1_76/A 8.58e-20
C16868 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# -5.42e-19
C16869 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# sky130_fd_sc_hd__conb_1_44/HI 1.37e-19
C16870 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 0.0179f
C16871 sky130_fd_sc_hd__inv_1_86/Y V_GND 0.136f
C16872 sky130_fd_sc_hd__dfbbn_1_2/a_581_47# V_GND 3.6e-19
C16873 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# RISING_COUNTER.COUNT_SUB_DFF12.Q 1.45e-21
C16874 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 0.00405f
C16875 sky130_fd_sc_hd__dfbbn_1_14/a_1159_47# sky130_fd_sc_hd__conb_1_18/HI -3.05e-20
C16876 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 5.84e-20
C16877 sky130_fd_sc_hd__dfbbn_1_38/a_1340_413# V_GND 2.23e-19
C16878 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# sky130_fd_sc_hd__conb_1_38/HI 0.00171f
C16879 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# V_LOW -0.00138f
C16880 sky130_fd_sc_hd__dfbbn_1_50/a_1340_413# V_GND 1.94e-19
C16881 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0.00614f
C16882 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 0.00271f
C16883 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 1.26e-19
C16884 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0173f
C16885 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# V_LOW -0.0109f
C16886 sky130_fd_sc_hd__conb_1_15/HI sky130_fd_sc_hd__dfbbn_1_15/a_1672_329# 2.44e-19
C16887 sky130_fd_sc_hd__nand2_1_5/a_113_47# V_LOW -1.78e-19
C16888 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# sky130_fd_sc_hd__conb_1_28/HI 0.00138f
C16889 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.432f
C16890 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_22/a_581_47# -7.91e-19
C16891 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# -0.0106f
C16892 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# sky130_fd_sc_hd__dfbbn_1_26/a_557_413# -0.0012f
C16893 sky130_fd_sc_hd__inv_1_71/A sky130_fd_sc_hd__inv_1_94/A 0.0395f
C16894 sky130_fd_sc_hd__dfbbn_1_9/a_1672_329# sky130_fd_sc_hd__conb_1_12/HI 4.53e-19
C16895 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 8.36e-20
C16896 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# sky130_fd_sc_hd__conb_1_21/HI 2.17e-20
C16897 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# -0.00282f
C16898 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 2.19e-20
C16899 sky130_fd_sc_hd__inv_1_111/Y sky130_fd_sc_hd__conb_1_34/HI 1.46e-20
C16900 sky130_fd_sc_hd__conb_1_24/LO sky130_fd_sc_hd__inv_16_0/Y 0.0186f
C16901 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# -5.33e-20
C16902 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# sky130_fd_sc_hd__dfbbn_1_31/a_557_413# -3.67e-20
C16903 sky130_fd_sc_hd__inv_1_63/Y V_LOW 0.111f
C16904 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# V_LOW -0.00389f
C16905 sky130_fd_sc_hd__dfbbn_1_27/a_557_413# V_GND 2.71e-19
C16906 sky130_fd_sc_hd__dfbbn_1_47/a_557_413# V_GND 1.87e-19
C16907 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__dfbbn_1_45/a_581_47# -2.6e-20
C16908 sky130_fd_sc_hd__dfbbn_1_11/a_1159_47# sky130_fd_sc_hd__conb_1_16/HI 0.00198f
C16909 sky130_fd_sc_hd__inv_1_95/A V_LOW 0.847f
C16910 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# RISING_COUNTER.COUNT_SUB_DFF5.Q 1.64e-20
C16911 sky130_fd_sc_hd__conb_1_23/HI sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 5.9e-19
C16912 sky130_fd_sc_hd__nand3_1_1/a_109_47# V_LOW -2.94e-19
C16913 RISING_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__inv_16_0/Y 0.0954f
C16914 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_647_21# -8.61e-20
C16915 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# sky130_fd_sc_hd__conb_1_17/HI 8.2e-21
C16916 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0.0485f
C16917 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# sky130_fd_sc_hd__conb_1_40/HI 0.0133f
C16918 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 2.72e-20
C16919 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 6.93e-21
C16920 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# V_LOW 0.00439f
C16921 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# sky130_fd_sc_hd__conb_1_25/HI 2.58e-19
C16922 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0166f
C16923 sky130_fd_sc_hd__dfbbn_1_0/a_1112_329# V_GND 7.43e-19
C16924 sky130_fd_sc_hd__dfbbn_1_31/a_891_329# FALLING_COUNTER.COUNT_SUB_DFF5.Q 1.93e-21
C16925 sky130_fd_sc_hd__dfbbn_1_38/a_1363_47# FALLING_COUNTER.COUNT_SUB_DFF12.Q 1.34e-19
C16926 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 6.57e-20
C16927 RISING_COUNTER.COUNT_SUB_DFF10.Q RISING_COUNTER.COUNT_SUB_DFF15.Q 1.73e-19
C16928 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0.00326f
C16929 sky130_fd_sc_hd__dfbbn_1_36/Q_N FALLING_COUNTER.COUNT_SUB_DFF13.Q 0.0163f
C16930 sky130_fd_sc_hd__inv_1_17/Y RISING_COUNTER.COUNT_SUB_DFF2.Q 1.48e-19
C16931 sky130_fd_sc_hd__dfbbn_1_7/a_1112_329# sky130_fd_sc_hd__inv_1_18/Y 0.00881f
C16932 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF6.Q 4.43e-21
C16933 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0043f
C16934 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# sky130_fd_sc_hd__dfbbn_1_18/a_581_47# -2.6e-20
C16935 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__inv_16_1/Y 0.0416f
C16936 sky130_fd_sc_hd__dfbbn_1_50/a_1672_329# FALLING_COUNTER.COUNT_SUB_DFF1.Q 0.00285f
C16937 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# V_GND 0.00228f
C16938 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# sky130_fd_sc_hd__dfbbn_1_44/a_941_21# -6.22e-19
C16939 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# -6.23e-21
C16940 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# sky130_fd_sc_hd__dfbbn_1_44/a_381_47# -0.00464f
C16941 sky130_fd_sc_hd__dfbbn_1_0/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF2.Q 5.12e-19
C16942 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# FULL_COUNTER.COUNT_SUB_DFF3.Q 0.00639f
C16943 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# sky130_fd_sc_hd__conb_1_32/HI 4.77e-19
C16944 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# FULL_COUNTER.COUNT_SUB_DFF10.Q 1.99e-20
C16945 sky130_fd_sc_hd__conb_1_4/HI FULL_COUNTER.COUNT_SUB_DFF3.Q 9.13e-21
C16946 sky130_fd_sc_hd__dfbbn_1_33/a_1340_413# sky130_fd_sc_hd__conb_1_35/HI 4.61e-19
C16947 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# RISING_COUNTER.COUNT_SUB_DFF3.Q 9.11e-20
C16948 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_941_21# -0.00171f
C16949 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# -3.72e-19
C16950 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# sky130_fd_sc_hd__inv_1_54/Y 4.43e-21
C16951 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# Reset 1.13e-19
C16952 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# sky130_fd_sc_hd__conb_1_40/HI 9.37e-21
C16953 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 4.43e-20
C16954 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# RISING_COUNTER.COUNT_SUB_DFF10.Q 0.0354f
C16955 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# sky130_fd_sc_hd__conb_1_27/LO 2.41e-20
C16956 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# sky130_fd_sc_hd__nand3_1_0/Y 2.54e-21
C16957 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00325f
C16958 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_58/Y 0.0717f
C16959 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# FALLING_COUNTER.COUNT_SUB_DFF3.Q 9.29e-19
C16960 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 6.92e-20
C16961 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__conb_1_35/HI 1.99e-19
C16962 sky130_fd_sc_hd__inv_16_2/Y sky130_fd_sc_hd__conb_1_12/HI 0.145f
C16963 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 2.35e-20
C16964 RISING_COUNTER.COUNT_SUB_DFF14.Q V_LOW 2.27f
C16965 sky130_fd_sc_hd__dfbbn_1_49/a_1159_47# sky130_fd_sc_hd__conb_1_38/HI -0.0024f
C16966 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# V_LOW 0.0035f
C16967 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# V_GND -0.005f
C16968 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 5.03e-19
C16969 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 4.19e-19
C16970 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 8.33e-19
C16971 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# FALLING_COUNTER.COUNT_SUB_DFF9.Q 0.0441f
C16972 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# V_LOW 0.00189f
C16973 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0.00517f
C16974 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__inv_1_22/Y 4.06e-21
C16975 sky130_fd_sc_hd__dfbbn_1_20/a_1340_413# RISING_COUNTER.COUNT_SUB_DFF11.Q 0.00113f
C16976 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# -5.42e-19
C16977 FALLING_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 3.28e-21
C16978 sky130_fd_sc_hd__conb_1_15/HI FULL_COUNTER.COUNT_SUB_DFF13.Q 0.0797f
C16979 sky130_fd_sc_hd__conb_1_15/LO V_LOW 0.151f
C16980 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 0.00165f
C16981 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 2.09e-21
C16982 sky130_fd_sc_hd__inv_1_94/Y sky130_fd_sc_hd__inv_1_68/A 4.7e-20
C16983 sky130_fd_sc_hd__nand3_1_0/a_193_47# V_LOW -4.71e-19
C16984 sky130_fd_sc_hd__conb_1_39/HI V_GND -0.089f
C16985 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# -1.67e-19
C16986 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# sky130_fd_sc_hd__dfbbn_1_32/a_381_47# -0.00565f
C16987 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# sky130_fd_sc_hd__dfbbn_1_32/a_941_21# -6.22e-19
C16988 FALLING_COUNTER.COUNT_SUB_DFF9.Q FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.664f
C16989 sky130_fd_sc_hd__conb_1_14/LO FULL_COUNTER.COUNT_SUB_DFF1.Q 0.00404f
C16990 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__inv_1_11/Y 0.117f
C16991 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 4.32e-19
C16992 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# sky130_fd_sc_hd__conb_1_22/LO 1.01e-19
C16993 FULL_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__conb_1_6/LO 0.00443f
C16994 sky130_fd_sc_hd__inv_1_72/Y sky130_fd_sc_hd__inv_1_76/A 0.0463f
C16995 sky130_fd_sc_hd__conb_1_18/HI sky130_fd_sc_hd__inv_16_2/Y 0.331f
C16996 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF13.Q 1.16e-19
C16997 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# sky130_fd_sc_hd__conb_1_48/HI -0.00117f
C16998 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# sky130_fd_sc_hd__inv_1_55/Y 0.00363f
C16999 FULL_COUNTER.COUNT_SUB_DFF0.Q sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0.203f
C17000 RISING_COUNTER.COUNT_SUB_DFF3.Q sky130_fd_sc_hd__inv_1_53/Y 9.85e-20
C17001 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# sky130_fd_sc_hd__conb_1_46/LO 0.0141f
C17002 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_57/Y 5.67e-20
C17003 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# V_LOW 0.0226f
C17004 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 2.01e-19
C17005 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# V_LOW 1.38e-19
C17006 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 1.51e-19
C17007 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 2.19e-19
C17008 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# sky130_fd_sc_hd__dfbbn_1_25/a_581_47# -7.91e-19
C17009 RISING_COUNTER.COUNT_SUB_DFF1.Q sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# 7.7e-19
C17010 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# sky130_fd_sc_hd__inv_1_57/Y 0.309f
C17011 sky130_fd_sc_hd__dfbbn_1_30/a_1159_47# sky130_fd_sc_hd__conb_1_40/HI 0.00125f
C17012 sky130_fd_sc_hd__inv_1_26/Y sky130_fd_sc_hd__inv_1_32/A 0.0443f
C17013 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_2/Y 0.0215f
C17014 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_31/Y 0.0113f
C17015 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# sky130_fd_sc_hd__inv_16_1/Y 0.0138f
C17016 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# sky130_fd_sc_hd__inv_1_56/Y 0.00265f
C17017 CLOCK_GEN.SR_Op.Q sky130_fd_sc_hd__nand2_1_0/Y 1.69e-19
C17018 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 1.31e-20
C17019 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 1.31e-20
C17020 sky130_fd_sc_hd__dfbbn_1_41/Q_N RISING_COUNTER.COUNT_SUB_DFF1.Q 0.0201f
C17021 sky130_fd_sc_hd__dfbbn_1_45/a_557_413# FALLING_COUNTER.COUNT_SUB_DFF8.Q 0.00226f
C17022 sky130_fd_sc_hd__dfbbn_1_25/a_1112_329# RISING_COUNTER.COUNT_SUB_DFF15.Q 0.00461f
C17023 FULL_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__inv_1_17/Y 0.0232f
C17024 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# FULL_COUNTER.COUNT_SUB_DFF7.Q 0.045f
C17025 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 0.00217f
C17026 sky130_fd_sc_hd__conb_1_28/HI V_GND -0.14f
C17027 FALLING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_36/a_1112_329# 1.1e-21
C17028 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# RISING_COUNTER.COUNT_SUB_DFF0.Q 6.76e-19
C17029 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# sky130_fd_sc_hd__inv_1_100/Y 3.71e-21
C17030 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# sky130_fd_sc_hd__inv_16_0/Y 0.00379f
C17031 sky130_fd_sc_hd__dfbbn_1_12/a_1672_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 2.3e-19
C17032 FULL_COUNTER.COUNT_SUB_DFF15.Q sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 0.166f
C17033 sky130_fd_sc_hd__dfbbn_1_33/a_557_413# V_GND 2.09e-19
C17034 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# FULL_COUNTER.COUNT_SUB_DFF15.Q 6.83e-20
C17035 sky130_fd_sc_hd__dfbbn_1_32/Q_N sky130_fd_sc_hd__inv_16_1/Y 0.0247f
C17036 sky130_fd_sc_hd__dfbbn_1_41/a_1112_329# V_GND 9.38e-19
C17037 sky130_fd_sc_hd__dfbbn_1_42/Q_N V_GND -0.00136f
C17038 sky130_fd_sc_hd__dfbbn_1_22/a_1159_47# sky130_fd_sc_hd__conb_1_32/HI -0.00236f
C17039 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# V_LOW 1.93e-19
C17040 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__dfbbn_1_25/a_381_47# 3.85e-19
C17041 sky130_fd_sc_hd__dfbbn_1_1/a_1112_329# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.02e-21
C17042 RISING_COUNTER.COUNT_SUB_DFF14.Q sky130_fd_sc_hd__dfbbn_1_20/a_27_47# 0.0321f
C17043 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# sky130_fd_sc_hd__inv_1_112/Y 2.83e-19
C17044 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF1.Q 0.0166f
C17045 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# -1.66e-19
C17046 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# sky130_fd_sc_hd__dfbbn_1_28/a_1672_329# -7.17e-20
C17047 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# sky130_fd_sc_hd__nand3_1_2/Y 0.0298f
C17048 sky130_fd_sc_hd__nand2_1_3/a_113_47# V_LOW -1.78e-19
C17049 sky130_fd_sc_hd__dfbbn_1_11/a_1363_47# FULL_COUNTER.COUNT_SUB_DFF1.Q 3.1e-19
C17050 sky130_fd_sc_hd__inv_1_75/Y sky130_fd_sc_hd__inv_1_67/Y 1.9e-19
C17051 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# -3.48e-20
C17052 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# sky130_fd_sc_hd__dfbbn_1_51/a_891_329# -2.2e-20
C17053 sky130_fd_sc_hd__inv_1_111/Y V_LOW 0.258f
C17054 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# sky130_fd_sc_hd__conb_1_35/HI 3.29e-20
C17055 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# Reset 0.00193f
C17056 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# Reset 6.81e-19
C17057 sky130_fd_sc_hd__nand2_8_6/a_27_47# RISING_COUNTER.COUNT_SUB_DFF4.Q 6.45e-20
C17058 sky130_fd_sc_hd__dfbbn_1_24/a_1112_329# V_GND 7.46e-19
C17059 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# CLOCK_GEN.SR_Op.Q 8.11e-21
C17060 sky130_fd_sc_hd__conb_1_7/HI sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 1.67e-21
C17061 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# sky130_fd_sc_hd__conb_1_34/HI 0.036f
C17062 sky130_fd_sc_hd__dfbbn_1_6/Q_N V_GND -0.00801f
C17063 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# FULL_COUNTER.COUNT_SUB_DFF1.Q 4.08e-19
C17064 sky130_fd_sc_hd__dfbbn_1_0/a_1159_47# sky130_fd_sc_hd__inv_1_7/Y 1.07e-19
C17065 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__inv_1_119/Y 1.2e-19
C17066 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__conb_1_5/LO 0.00147f
C17067 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# sky130_fd_sc_hd__conb_1_11/HI 3.18e-21
C17068 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# FULL_COUNTER.COUNT_SUB_DFF8.Q 0.00893f
C17069 sky130_fd_sc_hd__conb_1_3/LO sky130_fd_sc_hd__dfbbn_1_2/a_473_413# 0.00185f
C17070 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_16_1/Y 2.16e-21
C17071 sky130_fd_sc_hd__inv_1_43/A sky130_fd_sc_hd__inv_1_50/A 0.00663f
C17072 RISING_COUNTER.COUNT_SUB_DFF13.Q sky130_fd_sc_hd__inv_1_53/Y 0.0061f
C17073 sky130_fd_sc_hd__inv_1_110/Y sky130_fd_sc_hd__conb_1_44/HI 2.67e-19
C17074 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# -2.74e-21
C17075 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# sky130_fd_sc_hd__dfbbn_1_10/a_941_21# -7.6e-19
C17076 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# -0.00263f
C17077 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# RISING_COUNTER.COUNT_SUB_DFF2.Q 2.07e-20
C17078 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# CLOCK_GEN.SR_Op.Q 6.93e-20
C17079 sky130_fd_sc_hd__conb_1_9/HI sky130_fd_sc_hd__inv_16_2/Y 0.567f
C17080 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# sky130_fd_sc_hd__inv_16_1/Y 0.00159f
C17081 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# FULL_COUNTER.COUNT_SUB_DFF4.Q 0.00223f
C17082 sky130_fd_sc_hd__dfbbn_1_35/a_1363_47# RISING_COUNTER.COUNT_SUB_DFF7.Q 7.08e-20
C17083 sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 4.59e-19
C17084 sky130_fd_sc_hd__conb_1_4/HI FULL_COUNTER.COUNT_SUB_DFF5.Q 0.138f
C17085 sky130_fd_sc_hd__conb_1_1/LO FULL_COUNTER.COUNT_SUB_DFF3.Q 0.0013f
C17086 sky130_fd_sc_hd__conb_1_20/HI sky130_fd_sc_hd__inv_1_55/Y 6.06e-21
C17087 sky130_fd_sc_hd__conb_1_20/LO RISING_COUNTER.COUNT_SUB_DFF0.Q 1.21e-19
C17088 sky130_fd_sc_hd__conb_1_35/HI V_LOW 0.142f
C17089 sky130_fd_sc_hd__fill_4_69/VPB V_LOW 0.797f
C17090 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# sky130_fd_sc_hd__conb_1_51/HI 3.38e-19
C17091 sky130_fd_sc_hd__dfbbn_1_26/a_1672_329# sky130_fd_sc_hd__inv_1_55/Y 1.07e-21
C17092 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# sky130_fd_sc_hd__conb_1_5/LO 1.11e-20
C17093 FULL_COUNTER.COUNT_SUB_DFF12.Q sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 1.9e-19
C17094 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# sky130_fd_sc_hd__dfbbn_1_19/a_557_413# -0.0012f
C17095 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# -0.0026f
C17096 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# V_LOW 0.0101f
C17097 FULL_COUNTER.COUNT_SUB_DFF17.Q FULL_COUNTER.COUNT_SUB_DFF16.Q 0.043f
C17098 FALLING_COUNTER.COUNT_SUB_DFF6.Q sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# 6.71e-19
C17099 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# V_LOW 4.63e-19
C17100 sky130_fd_sc_hd__dfbbn_1_6/Q_N sky130_fd_sc_hd__inv_1_12/Y 0.0298f
C17101 V_LOW 0 0.948p
C17102 RISING_COUNTER.COUNT_SUB_DFF4.Q 0 1.57f
C17103 V_SENSE 0 35.5f
C17104 V_HIGH 0 22.3f
C17105 V_GND 0 0.434p
C17106 FULL_COUNTER.COUNT_SUB_DFF11.Q 0 0.951f
C17107 sky130_fd_sc_hd__conb_1_6/HI 0 0.446f
C17108 sky130_fd_sc_hd__inv_1_12/Y 0 0.196f
C17109 sky130_fd_sc_hd__inv_1_15/Y 0 0.274f
C17110 sky130_fd_sc_hd__inv_1_20/Y 0 0.233f
C17111 sky130_fd_sc_hd__conb_1_17/HI 0 0.562f
C17112 sky130_fd_sc_hd__inv_1_22/Y 0 0.197f
C17113 FULL_COUNTER.COUNT_SUB_DFF18.Q 0 1.16f
C17114 sky130_fd_sc_hd__conb_1_16/HI 0 0.467f
C17115 sky130_fd_sc_hd__conb_1_13/HI 0 0.518f
C17116 sky130_fd_sc_hd__inv_1_23/Y 0 0.163f
C17117 sky130_fd_sc_hd__conb_1_12/HI 0 0.458f
C17118 sky130_fd_sc_hd__inv_16_2/Y 0 5.89f
C17119 sky130_fd_sc_hd__inv_1_4/Y 0 0.246f
C17120 sky130_fd_sc_hd__inv_1_8/Y 0 0.24f
C17121 sky130_fd_sc_hd__conb_1_5/HI 0 0.514f
C17122 sky130_fd_sc_hd__conb_1_11/HI 0 0.468f
C17123 sky130_fd_sc_hd__inv_1_5/Y 0 0.22f
C17124 FULL_COUNTER.COUNT_SUB_DFF2.Q 0 1.18f
C17125 sky130_fd_sc_hd__conb_1_2/HI 0 0.53f
C17126 sky130_fd_sc_hd__inv_1_9/Y 0 0.175f
C17127 sky130_fd_sc_hd__conb_1_0/HI 0 0.481f
C17128 sky130_fd_sc_hd__inv_1_10/Y 0 0.232f
C17129 sky130_fd_sc_hd__conb_1_21/HI 0 0.5f
C17130 sky130_fd_sc_hd__inv_1_53/Y 0 0.19f
C17131 sky130_fd_sc_hd__conb_1_22/HI 0 0.486f
C17132 RISING_COUNTER.COUNT_SUB_DFF15.Q 0 0.572f
C17133 sky130_fd_sc_hd__conb_1_26/HI 0 0.428f
C17134 sky130_fd_sc_hd__inv_1_57/Y 0 0.174f
C17135 sky130_fd_sc_hd__inv_1_58/Y 0 0.173f
C17136 sky130_fd_sc_hd__inv_1_112/Y 0 0.226f
C17137 sky130_fd_sc_hd__conb_1_30/HI 0 0.559f
C17138 sky130_fd_sc_hd__conb_1_28/HI 0 0.498f
C17139 sky130_fd_sc_hd__inv_1_60/Y 0 0.2f
C17140 RISING_COUNTER.COUNT_SUB_DFF6.Q 0 1.46f
C17141 sky130_fd_sc_hd__conb_1_24/HI 0 0.51f
C17142 RISING_COUNTER.COUNT_SUB_DFF3.Q 0 1.14f
C17143 sky130_fd_sc_hd__inv_1_63/Y 0 0.727f
C17144 sky130_fd_sc_hd__nand2_8_9/Y 0 0.702f
C17145 sky130_fd_sc_hd__inv_1_65/Y 0 0.265f
C17146 sky130_fd_sc_hd__inv_1_59/Y 0 0.201f
C17147 RISING_COUNTER.COUNT_SUB_DFF5.Q 0 1.24f
C17148 sky130_fd_sc_hd__inv_1_90/Y 0 0.231f
C17149 sky130_fd_sc_hd__nand3_1_1/Y 0 0.304f
C17150 sky130_fd_sc_hd__inv_1_93/A 0 0.915f
C17151 sky130_fd_sc_hd__inv_1_70/A 0 0.86f
C17152 sky130_fd_sc_hd__inv_1_68/A 0 0.904f
C17153 sky130_fd_sc_hd__inv_1_86/Y 0 0.218f
C17154 sky130_fd_sc_hd__inv_1_97/Y 0 0.196f
C17155 sky130_fd_sc_hd__inv_1_80/A 0 0.567f
C17156 sky130_fd_sc_hd__nand2_1_0/Y 0 0.221f
C17157 sky130_fd_sc_hd__inv_2_0/Y 0 2.28f
C17158 sky130_fd_sc_hd__inv_1_78/A 0 0.25f
C17159 sky130_fd_sc_hd__nand2_8_2/A 0 0.717f
C17160 sky130_fd_sc_hd__inv_1_75/A 0 0.745f
C17161 sky130_fd_sc_hd__inv_1_76/A 0 3.69f
C17162 sky130_fd_sc_hd__inv_1_67/Y 0 0.917f
C17163 sky130_fd_sc_hd__inv_1_45/A 0 0.365f
C17164 sky130_fd_sc_hd__nand2_8_3/Y 0 0.744f
C17165 sky130_fd_sc_hd__nand3_1_2/B 0 0.806f
C17166 sky130_fd_sc_hd__inv_1_97/A 0 0.251f
C17167 sky130_fd_sc_hd__inv_1_105/Y 0 0.214f
C17168 sky130_fd_sc_hd__conb_1_45/HI 0 0.433f
C17169 sky130_fd_sc_hd__conb_1_46/HI 0 0.442f
C17170 sky130_fd_sc_hd__inv_1_108/Y 0 0.348f
C17171 sky130_fd_sc_hd__inv_1_106/Y 0 0.156f
C17172 FALLING_COUNTER.COUNT_SUB_DFF8.Q 0 1.65f
C17173 sky130_fd_sc_hd__inv_1_99/Y 0 0.199f
C17174 sky130_fd_sc_hd__inv_16_1/Y 0 3.71f
C17175 sky130_fd_sc_hd__conb_1_35/HI 0 0.464f
C17176 sky130_fd_sc_hd__inv_1_101/Y 0 0.161f
C17177 sky130_fd_sc_hd__inv_1_100/Y 0 0.189f
C17178 sky130_fd_sc_hd__conb_1_41/HI 0 0.455f
C17179 sky130_fd_sc_hd__inv_1_50/Y 0 0.226f
C17180 sky130_fd_sc_hd__inv_1_50/A 0 1.02f
C17181 sky130_fd_sc_hd__inv_1_43/A 0 0.265f
C17182 sky130_fd_sc_hd__conb_1_40/HI 0 0.506f
C17183 FALLING_COUNTER.COUNT_SUB_DFF0.Q 0 2.37f
C17184 sky130_fd_sc_hd__inv_1_47/Y 0 0.282f
C17185 sky130_fd_sc_hd__inv_1_3/Y 0 0.162f
C17186 sky130_fd_sc_hd__inv_1_2/A 0 0.164f
C17187 sky130_fd_sc_hd__inv_1_2/Y 0 0.183f
C17188 sky130_fd_sc_hd__inv_1_31/Y 0 0.163f
C17189 sky130_fd_sc_hd__inv_1_31/A 0 0.161f
C17190 sky130_fd_sc_hd__inv_1_1/Y 0 0.171f
C17191 sky130_fd_sc_hd__inv_1_34/A 0 0.162f
C17192 sky130_fd_sc_hd__inv_1_32/Y 0 0.16f
C17193 sky130_fd_sc_hd__inv_1_32/A 0 0.16f
C17194 sky130_fd_sc_hd__inv_1_26/Y 0 0.161f
C17195 sky130_fd_sc_hd__inv_1_27/Y 0 0.17f
C17196 sky130_fd_sc_hd__inv_1_28/Y 0 0.162f
C17197 sky130_fd_sc_hd__inv_1_33/Y 0 0.165f
C17198 sky130_fd_sc_hd__inv_1_0/A 0 0.205f
C17199 sky130_fd_sc_hd__inv_1_3/A 0 0.267f
C17200 FULL_COUNTER.COUNT_SUB_DFF10.Q 0 1.26f
C17201 FULL_COUNTER.COUNT_SUB_DFF9.Q 0 1.03f
C17202 sky130_fd_sc_hd__inv_1_11/Y 0 0.171f
C17203 FULL_COUNTER.COUNT_SUB_DFF8.Q 0 1.16f
C17204 FULL_COUNTER.COUNT_SUB_DFF5.Q 0 1.32f
C17205 sky130_fd_sc_hd__inv_1_13/Y 0 0.141f
C17206 FULL_COUNTER.COUNT_SUB_DFF4.Q 0 2.02f
C17207 FULL_COUNTER.COUNT_SUB_DFF13.Q 0 1.58f
C17208 sky130_fd_sc_hd__inv_1_18/Y 0 0.285f
C17209 FULL_COUNTER.COUNT_SUB_DFF1.Q 0 0.936f
C17210 FULL_COUNTER.COUNT_SUB_DFF16.Q 0 0.778f
C17211 sky130_fd_sc_hd__inv_1_19/Y 0 0.217f
C17212 transmission_gate_0/GN 0 0.099f
C17213 sky130_fd_sc_hd__inv_2_0/A 0 0.25f
C17214 sky130_fd_sc_hd__inv_1_119/Y 0 0.926f
C17215 sky130_fd_sc_hd__inv_1_72/A 0 0.272f
C17216 RISING_COUNTER.COUNT_SUB_DFF13.Q 0 0.968f
C17217 Reset 0 6.76f
C17218 sky130_fd_sc_hd__nor2_1_0/Y 0 0.135f
C17219 RISING_COUNTER.COUNT_SUB_DFF2.Q 0 0.989f
C17220 sky130_fd_sc_hd__inv_16_0/Y 0 5.2f
C17221 sky130_fd_sc_hd__nand3_1_0/Y 0 0.826f
C17222 CLOCK_GEN.SR_Op.Q 0 1.48f
C17223 sky130_fd_sc_hd__inv_1_56/Y 0 0.145f
C17224 RISING_COUNTER.COUNT_SUB_DFF11.Q 0 0.929f
C17225 RISING_COUNTER.COUNT_SUB_DFF0.Q 0 1.73f
C17226 sky130_fd_sc_hd__inv_1_70/Y 0 0.22f
C17227 sky130_fd_sc_hd__inv_1_66/Y 0 0.777f
C17228 sky130_fd_sc_hd__inv_1_71/Y 0 0.35f
C17229 sky130_fd_sc_hd__inv_1_55/Y 0 0.2f
C17230 sky130_fd_sc_hd__inv_1_94/A 0 0.811f
C17231 sky130_fd_sc_hd__inv_1_40/A 0 0.157f
C17232 sky130_fd_sc_hd__inv_1_44/A 0 0.169f
C17233 sky130_fd_sc_hd__inv_1_39/A 0 0.199f
C17234 sky130_fd_sc_hd__conb_1_32/HI 0 0.534f
C17235 sky130_fd_sc_hd__inv_1_61/Y 0 0.235f
C17236 sky130_fd_sc_hd__inv_1_95/A 0 0.719f
C17237 sky130_fd_sc_hd__conb_1_31/HI 0 0.444f
C17238 RISING_COUNTER.COUNT_SUB_DFF9.Q 0 1.76f
C17239 sky130_fd_sc_hd__inv_1_62/Y 0 0.145f
C17240 sky130_fd_sc_hd__inv_1_83/Y 0 0.298f
C17241 sky130_fd_sc_hd__inv_1_85/Y 0 0.229f
C17242 RISING_COUNTER.COUNT_SUB_DFF7.Q 0 0.76f
C17243 sky130_fd_sc_hd__inv_1_95/Y 0 0.192f
C17244 sky130_fd_sc_hd__inv_1_75/Y 0 0.658f
C17245 sky130_fd_sc_hd__inv_1_42/Y 0 0.154f
C17246 sky130_fd_sc_hd__inv_1_43/Y 0 0.156f
C17247 sky130_fd_sc_hd__inv_1_85/A 0 0.249f
C17248 sky130_fd_sc_hd__inv_1_74/Y 0 0.28f
C17249 sky130_fd_sc_hd__inv_1_92/Y 0 0.342f
C17250 sky130_fd_sc_hd__inv_1_91/A 0 0.173f
C17251 sky130_fd_sc_hd__inv_1_91/Y 0 0.23f
C17252 sky130_fd_sc_hd__inv_1_103/Y 0 0.237f
C17253 sky130_fd_sc_hd__inv_1_107/Y 0 0.189f
C17254 FALLING_COUNTER.COUNT_SUB_DFF13.Q 0 0.956f
C17255 FALLING_COUNTER.COUNT_SUB_DFF9.Q 0 1.54f
C17256 FALLING_COUNTER.COUNT_SUB_DFF11.Q 0 1.23f
C17257 FALLING_COUNTER.COUNT_SUB_DFF10.Q 0 2.27f
C17258 sky130_fd_sc_hd__conb_1_44/HI 0 0.442f
C17259 FALLING_COUNTER.COUNT_SUB_DFF5.Q 0 1.24f
C17260 sky130_fd_sc_hd__conb_1_47/HI 0 0.456f
C17261 sky130_fd_sc_hd__inv_1_6/Y 0 0.171f
C17262 FULL_COUNTER.COUNT_SUB_DFF7.Q 0 1.87f
C17263 sky130_fd_sc_hd__fill_4_73/VPB 0 4.66f
C17264 sky130_fd_sc_hd__dfbbn_1_5/Q_N 0 0.0135f
C17265 sky130_fd_sc_hd__dfbbn_1_5/a_1555_47# 0 0.00871f
C17266 sky130_fd_sc_hd__dfbbn_1_5/a_2136_47# 0 0.133f
C17267 sky130_fd_sc_hd__dfbbn_1_5/a_791_47# 0 0.0125f
C17268 sky130_fd_sc_hd__dfbbn_1_5/a_381_47# 0 0.0218f
C17269 sky130_fd_sc_hd__dfbbn_1_5/a_1256_413# 0 0.12f
C17270 sky130_fd_sc_hd__dfbbn_1_5/a_1415_315# 0 0.394f
C17271 sky130_fd_sc_hd__dfbbn_1_5/a_941_21# 0 0.245f
C17272 sky130_fd_sc_hd__dfbbn_1_5/a_473_413# 0 0.119f
C17273 sky130_fd_sc_hd__dfbbn_1_5/a_647_21# 0 0.24f
C17274 sky130_fd_sc_hd__dfbbn_1_5/a_193_47# 0 0.27f
C17275 sky130_fd_sc_hd__dfbbn_1_5/a_27_47# 0 0.492f
C17276 sky130_fd_sc_hd__nand2_8_1/a_27_47# 0 0.083f
C17277 sky130_fd_sc_hd__conb_1_18/HI 0 0.461f
C17278 sky130_fd_sc_hd__inv_1_54/Y 0 0.196f
C17279 sky130_fd_sc_hd__inv_1_68/Y 0 0.0961f
C17280 sky130_fd_sc_hd__conb_1_49/HI 0 0.443f
C17281 sky130_fd_sc_hd__dfbbn_1_4/Q_N 0 0.0135f
C17282 sky130_fd_sc_hd__dfbbn_1_4/a_1555_47# 0 0.00871f
C17283 sky130_fd_sc_hd__dfbbn_1_4/a_2136_47# 0 0.133f
C17284 sky130_fd_sc_hd__dfbbn_1_4/a_791_47# 0 0.0125f
C17285 sky130_fd_sc_hd__dfbbn_1_4/a_381_47# 0 0.0218f
C17286 sky130_fd_sc_hd__dfbbn_1_4/a_1256_413# 0 0.12f
C17287 sky130_fd_sc_hd__dfbbn_1_4/a_1415_315# 0 0.394f
C17288 sky130_fd_sc_hd__dfbbn_1_4/a_941_21# 0 0.245f
C17289 sky130_fd_sc_hd__dfbbn_1_4/a_473_413# 0 0.119f
C17290 sky130_fd_sc_hd__dfbbn_1_4/a_647_21# 0 0.24f
C17291 sky130_fd_sc_hd__dfbbn_1_4/a_193_47# 0 0.27f
C17292 sky130_fd_sc_hd__dfbbn_1_4/a_27_47# 0 0.492f
C17293 sky130_fd_sc_hd__conb_1_34/HI 0 0.482f
C17294 sky130_fd_sc_hd__nand2_8_0/a_27_47# 0 0.083f
C17295 sky130_fd_sc_hd__conb_1_9/LO 0 0.166f
C17296 FULL_COUNTER.COUNT_SUB_DFF3.Q 0 1f
C17297 sky130_fd_sc_hd__inv_1_79/A 0 0.153f
C17298 sky130_fd_sc_hd__dfbbn_1_3/Q_N 0 0.0135f
C17299 sky130_fd_sc_hd__dfbbn_1_3/a_1555_47# 0 0.00871f
C17300 sky130_fd_sc_hd__dfbbn_1_3/a_2136_47# 0 0.133f
C17301 sky130_fd_sc_hd__dfbbn_1_3/a_791_47# 0 0.0125f
C17302 sky130_fd_sc_hd__dfbbn_1_3/a_381_47# 0 0.0218f
C17303 sky130_fd_sc_hd__dfbbn_1_3/a_1256_413# 0 0.12f
C17304 sky130_fd_sc_hd__dfbbn_1_3/a_1415_315# 0 0.394f
C17305 sky130_fd_sc_hd__dfbbn_1_3/a_941_21# 0 0.245f
C17306 sky130_fd_sc_hd__dfbbn_1_3/a_473_413# 0 0.119f
C17307 sky130_fd_sc_hd__dfbbn_1_3/a_647_21# 0 0.24f
C17308 sky130_fd_sc_hd__dfbbn_1_3/a_193_47# 0 0.27f
C17309 sky130_fd_sc_hd__dfbbn_1_3/a_27_47# 0 0.492f
C17310 sky130_fd_sc_hd__conb_1_37/HI 0 0.461f
C17311 sky130_fd_sc_hd__conb_1_8/LO 0 0.166f
C17312 sky130_fd_sc_hd__conb_1_33/HI 0 0.445f
C17313 sky130_fd_sc_hd__dfbbn_1_2/Q_N 0 0.0135f
C17314 sky130_fd_sc_hd__dfbbn_1_2/a_1555_47# 0 0.00871f
C17315 sky130_fd_sc_hd__dfbbn_1_2/a_2136_47# 0 0.133f
C17316 sky130_fd_sc_hd__dfbbn_1_2/a_791_47# 0 0.0125f
C17317 sky130_fd_sc_hd__dfbbn_1_2/a_381_47# 0 0.0218f
C17318 sky130_fd_sc_hd__dfbbn_1_2/a_1256_413# 0 0.12f
C17319 sky130_fd_sc_hd__dfbbn_1_2/a_1415_315# 0 0.394f
C17320 sky130_fd_sc_hd__dfbbn_1_2/a_941_21# 0 0.245f
C17321 sky130_fd_sc_hd__dfbbn_1_2/a_473_413# 0 0.119f
C17322 sky130_fd_sc_hd__dfbbn_1_2/a_647_21# 0 0.24f
C17323 sky130_fd_sc_hd__dfbbn_1_2/a_193_47# 0 0.27f
C17324 sky130_fd_sc_hd__dfbbn_1_2/a_27_47# 0 0.492f
C17325 sky130_fd_sc_hd__conb_1_7/LO 0 0.166f
C17326 sky130_fd_sc_hd__dfbbn_1_1/Q_N 0 0.0135f
C17327 sky130_fd_sc_hd__dfbbn_1_1/a_1555_47# 0 0.00871f
C17328 sky130_fd_sc_hd__dfbbn_1_1/a_2136_47# 0 0.133f
C17329 sky130_fd_sc_hd__dfbbn_1_1/a_791_47# 0 0.0125f
C17330 sky130_fd_sc_hd__dfbbn_1_1/a_381_47# 0 0.0218f
C17331 sky130_fd_sc_hd__dfbbn_1_1/a_1256_413# 0 0.12f
C17332 sky130_fd_sc_hd__dfbbn_1_1/a_1415_315# 0 0.394f
C17333 sky130_fd_sc_hd__dfbbn_1_1/a_941_21# 0 0.245f
C17334 sky130_fd_sc_hd__dfbbn_1_1/a_473_413# 0 0.119f
C17335 sky130_fd_sc_hd__dfbbn_1_1/a_647_21# 0 0.24f
C17336 sky130_fd_sc_hd__dfbbn_1_1/a_193_47# 0 0.27f
C17337 sky130_fd_sc_hd__dfbbn_1_1/a_27_47# 0 0.492f
C17338 sky130_fd_sc_hd__conb_1_6/LO 0 0.166f
C17339 sky130_fd_sc_hd__inv_1_109/Y 0 0.149f
C17340 sky130_fd_sc_hd__inv_1_88/Y 0 0.188f
C17341 sky130_fd_sc_hd__dfbbn_1_0/Q_N 0 0.0135f
C17342 sky130_fd_sc_hd__dfbbn_1_0/a_1555_47# 0 0.00871f
C17343 sky130_fd_sc_hd__dfbbn_1_0/a_2136_47# 0 0.133f
C17344 sky130_fd_sc_hd__dfbbn_1_0/a_791_47# 0 0.0125f
C17345 sky130_fd_sc_hd__dfbbn_1_0/a_381_47# 0 0.0218f
C17346 sky130_fd_sc_hd__dfbbn_1_0/a_1256_413# 0 0.12f
C17347 sky130_fd_sc_hd__dfbbn_1_0/a_1415_315# 0 0.394f
C17348 sky130_fd_sc_hd__dfbbn_1_0/a_941_21# 0 0.245f
C17349 sky130_fd_sc_hd__dfbbn_1_0/a_473_413# 0 0.119f
C17350 sky130_fd_sc_hd__dfbbn_1_0/a_647_21# 0 0.24f
C17351 sky130_fd_sc_hd__dfbbn_1_0/a_193_47# 0 0.27f
C17352 sky130_fd_sc_hd__dfbbn_1_0/a_27_47# 0 0.492f
C17353 sky130_fd_sc_hd__nand2_1_3/Y 0 0.0557f
C17354 sky130_fd_sc_hd__conb_1_5/LO 0 0.166f
C17355 sky130_fd_sc_hd__conb_1_8/HI 0 0.449f
C17356 FALLING_COUNTER.COUNT_SUB_DFF1.Q 0 1.27f
C17357 sky130_fd_sc_hd__conb_1_4/LO 0 0.166f
C17358 sky130_fd_sc_hd__inv_1_51/Y 0 0.0961f
C17359 sky130_fd_sc_hd__conb_1_42/HI 0 0.44f
C17360 sky130_fd_sc_hd__inv_1_21/Y 0 0.209f
C17361 RISING_COUNTER.COUNT_SUB_DFF10.Q 0 1.73f
C17362 sky130_fd_sc_hd__conb_1_3/LO 0 0.166f
C17363 sky130_fd_sc_hd__nand3_1_2/Y 0 0.406f
C17364 sky130_fd_sc_hd__inv_1_102/Y 0 0.277f
C17365 sky130_fd_sc_hd__conb_1_19/LO 0 0.166f
C17366 sky130_fd_sc_hd__conb_1_2/LO 0 0.166f
C17367 sky130_fd_sc_hd__inv_1_93/Y 0 0.0961f
C17368 sky130_fd_sc_hd__inv_1_51/A 0 0.852f
C17369 sky130_fd_sc_hd__conb_1_18/LO 0 0.166f
C17370 sky130_fd_sc_hd__conb_1_29/LO 0 0.166f
C17371 sky130_fd_sc_hd__conb_1_1/LO 0 0.166f
C17372 sky130_fd_sc_hd__conb_1_17/LO 0 0.166f
C17373 sky130_fd_sc_hd__conb_1_28/LO 0 0.166f
C17374 sky130_fd_sc_hd__conb_1_39/LO 0 0.166f
C17375 sky130_fd_sc_hd__inv_1_72/Y 0 0.154f
C17376 sky130_fd_sc_hd__conb_1_0/LO 0 0.166f
C17377 sky130_fd_sc_hd__conb_1_9/HI 0 0.458f
C17378 sky130_fd_sc_hd__conb_1_38/HI 0 0.533f
C17379 sky130_fd_sc_hd__conb_1_49/LO 0 0.166f
C17380 sky130_fd_sc_hd__conb_1_16/LO 0 0.166f
C17381 sky130_fd_sc_hd__conb_1_27/LO 0 0.166f
C17382 sky130_fd_sc_hd__conb_1_38/LO 0 0.166f
C17383 sky130_fd_sc_hd__inv_1_16/Y 0 0.164f
C17384 sky130_fd_sc_hd__conb_1_15/LO 0 0.166f
C17385 sky130_fd_sc_hd__conb_1_26/LO 0 0.166f
C17386 sky130_fd_sc_hd__conb_1_37/LO 0 0.166f
C17387 sky130_fd_sc_hd__conb_1_48/LO 0 0.166f
C17388 sky130_fd_sc_hd__conb_1_27/HI 0 0.474f
C17389 sky130_fd_sc_hd__inv_1_69/Y 0 0.295f
C17390 sky130_fd_sc_hd__conb_1_14/LO 0 0.166f
C17391 sky130_fd_sc_hd__conb_1_25/LO 0 0.166f
C17392 sky130_fd_sc_hd__conb_1_36/LO 0 0.166f
C17393 sky130_fd_sc_hd__conb_1_47/LO 0 0.166f
C17394 sky130_fd_sc_hd__conb_1_3/HI 0 0.477f
C17395 sky130_fd_sc_hd__dfbbn_1_19/Q_N 0 0.0135f
C17396 sky130_fd_sc_hd__dfbbn_1_19/a_1555_47# 0 0.00871f
C17397 sky130_fd_sc_hd__dfbbn_1_19/a_2136_47# 0 0.133f
C17398 sky130_fd_sc_hd__dfbbn_1_19/a_791_47# 0 0.0125f
C17399 sky130_fd_sc_hd__dfbbn_1_19/a_381_47# 0 0.0218f
C17400 sky130_fd_sc_hd__dfbbn_1_19/a_1256_413# 0 0.12f
C17401 sky130_fd_sc_hd__dfbbn_1_19/a_1415_315# 0 0.394f
C17402 sky130_fd_sc_hd__dfbbn_1_19/a_941_21# 0 0.245f
C17403 sky130_fd_sc_hd__dfbbn_1_19/a_473_413# 0 0.119f
C17404 sky130_fd_sc_hd__dfbbn_1_19/a_647_21# 0 0.24f
C17405 sky130_fd_sc_hd__dfbbn_1_19/a_193_47# 0 0.27f
C17406 sky130_fd_sc_hd__dfbbn_1_19/a_27_47# 0 0.492f
C17407 sky130_fd_sc_hd__conb_1_39/HI 0 0.453f
C17408 sky130_fd_sc_hd__conb_1_13/LO 0 0.166f
C17409 sky130_fd_sc_hd__conb_1_24/LO 0 0.166f
C17410 sky130_fd_sc_hd__conb_1_46/LO 0 0.166f
C17411 sky130_fd_sc_hd__conb_1_35/LO 0 0.166f
C17412 sky130_fd_sc_hd__dfbbn_1_18/Q_N 0 0.0135f
C17413 sky130_fd_sc_hd__dfbbn_1_18/a_1555_47# 0 0.00871f
C17414 sky130_fd_sc_hd__dfbbn_1_18/a_2136_47# 0 0.133f
C17415 sky130_fd_sc_hd__dfbbn_1_18/a_791_47# 0 0.0125f
C17416 sky130_fd_sc_hd__dfbbn_1_18/a_381_47# 0 0.0218f
C17417 sky130_fd_sc_hd__dfbbn_1_18/a_1256_413# 0 0.12f
C17418 sky130_fd_sc_hd__dfbbn_1_18/a_1415_315# 0 0.394f
C17419 sky130_fd_sc_hd__dfbbn_1_18/a_941_21# 0 0.245f
C17420 sky130_fd_sc_hd__dfbbn_1_18/a_473_413# 0 0.119f
C17421 sky130_fd_sc_hd__dfbbn_1_18/a_647_21# 0 0.24f
C17422 sky130_fd_sc_hd__dfbbn_1_18/a_193_47# 0 0.27f
C17423 sky130_fd_sc_hd__dfbbn_1_18/a_27_47# 0 0.492f
C17424 sky130_fd_sc_hd__dfbbn_1_29/Q_N 0 0.0135f
C17425 sky130_fd_sc_hd__dfbbn_1_29/a_1555_47# 0 0.00871f
C17426 sky130_fd_sc_hd__dfbbn_1_29/a_2136_47# 0 0.133f
C17427 sky130_fd_sc_hd__dfbbn_1_29/a_791_47# 0 0.0125f
C17428 sky130_fd_sc_hd__dfbbn_1_29/a_381_47# 0 0.0218f
C17429 sky130_fd_sc_hd__dfbbn_1_29/a_1256_413# 0 0.12f
C17430 sky130_fd_sc_hd__dfbbn_1_29/a_1415_315# 0 0.394f
C17431 sky130_fd_sc_hd__dfbbn_1_29/a_941_21# 0 0.245f
C17432 sky130_fd_sc_hd__dfbbn_1_29/a_473_413# 0 0.119f
C17433 sky130_fd_sc_hd__dfbbn_1_29/a_647_21# 0 0.24f
C17434 sky130_fd_sc_hd__dfbbn_1_29/a_193_47# 0 0.27f
C17435 sky130_fd_sc_hd__dfbbn_1_29/a_27_47# 0 0.492f
C17436 sky130_fd_sc_hd__inv_1_71/A 0 1.46f
C17437 sky130_fd_sc_hd__fill_4_84/VPB 0 4.66f
C17438 sky130_fd_sc_hd__conb_1_51/HI 0 0.483f
C17439 sky130_fd_sc_hd__conb_1_12/LO 0 0.166f
C17440 sky130_fd_sc_hd__conb_1_23/LO 0 0.166f
C17441 sky130_fd_sc_hd__inv_1_64/A 0 0.9f
C17442 sky130_fd_sc_hd__conb_1_34/LO 0 0.166f
C17443 sky130_fd_sc_hd__conb_1_45/LO 0 0.166f
C17444 sky130_fd_sc_hd__dfbbn_1_17/Q_N 0 0.0135f
C17445 sky130_fd_sc_hd__dfbbn_1_17/a_1555_47# 0 0.00871f
C17446 sky130_fd_sc_hd__dfbbn_1_17/a_2136_47# 0 0.133f
C17447 sky130_fd_sc_hd__dfbbn_1_17/a_791_47# 0 0.0125f
C17448 sky130_fd_sc_hd__dfbbn_1_17/a_381_47# 0 0.0218f
C17449 sky130_fd_sc_hd__dfbbn_1_17/a_1256_413# 0 0.12f
C17450 sky130_fd_sc_hd__dfbbn_1_17/a_1415_315# 0 0.394f
C17451 sky130_fd_sc_hd__dfbbn_1_17/a_941_21# 0 0.245f
C17452 sky130_fd_sc_hd__dfbbn_1_17/a_473_413# 0 0.119f
C17453 sky130_fd_sc_hd__dfbbn_1_17/a_647_21# 0 0.24f
C17454 sky130_fd_sc_hd__dfbbn_1_17/a_193_47# 0 0.27f
C17455 sky130_fd_sc_hd__dfbbn_1_17/a_27_47# 0 0.492f
C17456 sky130_fd_sc_hd__dfbbn_1_28/Q_N 0 0.0135f
C17457 sky130_fd_sc_hd__dfbbn_1_28/a_1555_47# 0 0.00871f
C17458 sky130_fd_sc_hd__dfbbn_1_28/a_2136_47# 0 0.133f
C17459 sky130_fd_sc_hd__dfbbn_1_28/a_791_47# 0 0.0125f
C17460 sky130_fd_sc_hd__dfbbn_1_28/a_381_47# 0 0.0218f
C17461 sky130_fd_sc_hd__dfbbn_1_28/a_1256_413# 0 0.12f
C17462 sky130_fd_sc_hd__dfbbn_1_28/a_1415_315# 0 0.394f
C17463 sky130_fd_sc_hd__dfbbn_1_28/a_941_21# 0 0.245f
C17464 sky130_fd_sc_hd__dfbbn_1_28/a_473_413# 0 0.119f
C17465 sky130_fd_sc_hd__dfbbn_1_28/a_647_21# 0 0.24f
C17466 sky130_fd_sc_hd__dfbbn_1_28/a_193_47# 0 0.27f
C17467 sky130_fd_sc_hd__dfbbn_1_28/a_27_47# 0 0.492f
C17468 sky130_fd_sc_hd__dfbbn_1_39/Q_N 0 0.0135f
C17469 sky130_fd_sc_hd__dfbbn_1_39/a_1555_47# 0 0.00871f
C17470 sky130_fd_sc_hd__dfbbn_1_39/a_2136_47# 0 0.133f
C17471 sky130_fd_sc_hd__dfbbn_1_39/a_791_47# 0 0.0125f
C17472 sky130_fd_sc_hd__dfbbn_1_39/a_381_47# 0 0.0218f
C17473 sky130_fd_sc_hd__dfbbn_1_39/a_1256_413# 0 0.12f
C17474 sky130_fd_sc_hd__dfbbn_1_39/a_1415_315# 0 0.394f
C17475 sky130_fd_sc_hd__dfbbn_1_39/a_941_21# 0 0.245f
C17476 sky130_fd_sc_hd__dfbbn_1_39/a_473_413# 0 0.119f
C17477 sky130_fd_sc_hd__dfbbn_1_39/a_647_21# 0 0.24f
C17478 sky130_fd_sc_hd__dfbbn_1_39/a_193_47# 0 0.27f
C17479 sky130_fd_sc_hd__dfbbn_1_39/a_27_47# 0 0.492f
C17480 FALLING_COUNTER.COUNT_SUB_DFF12.Q 0 0.903f
C17481 sky130_fd_sc_hd__inv_1_98/Y 0 0.189f
C17482 FALLING_COUNTER.COUNT_SUB_DFF7.Q 0 1.77f
C17483 sky130_fd_sc_hd__conb_1_33/LO 0 0.166f
C17484 sky130_fd_sc_hd__conb_1_44/LO 0 0.166f
C17485 sky130_fd_sc_hd__conb_1_11/LO 0 0.166f
C17486 sky130_fd_sc_hd__conb_1_22/LO 0 0.166f
C17487 RISING_COUNTER.COUNT_SUB_DFF12.Q 0 1.96f
C17488 sky130_fd_sc_hd__conb_1_4/HI 0 0.493f
C17489 sky130_fd_sc_hd__dfbbn_1_16/Q_N 0 0.0135f
C17490 sky130_fd_sc_hd__dfbbn_1_16/a_1555_47# 0 0.00871f
C17491 sky130_fd_sc_hd__dfbbn_1_16/a_2136_47# 0 0.133f
C17492 sky130_fd_sc_hd__dfbbn_1_16/a_791_47# 0 0.0125f
C17493 sky130_fd_sc_hd__dfbbn_1_16/a_381_47# 0 0.0218f
C17494 sky130_fd_sc_hd__dfbbn_1_16/a_1256_413# 0 0.12f
C17495 sky130_fd_sc_hd__dfbbn_1_16/a_1415_315# 0 0.394f
C17496 sky130_fd_sc_hd__dfbbn_1_16/a_941_21# 0 0.245f
C17497 sky130_fd_sc_hd__dfbbn_1_16/a_473_413# 0 0.119f
C17498 sky130_fd_sc_hd__dfbbn_1_16/a_647_21# 0 0.24f
C17499 sky130_fd_sc_hd__dfbbn_1_16/a_193_47# 0 0.27f
C17500 sky130_fd_sc_hd__dfbbn_1_16/a_27_47# 0 0.492f
C17501 sky130_fd_sc_hd__dfbbn_1_27/Q_N 0 0.0135f
C17502 sky130_fd_sc_hd__conb_1_23/HI 0 0.414f
C17503 sky130_fd_sc_hd__dfbbn_1_27/a_1555_47# 0 0.00871f
C17504 sky130_fd_sc_hd__dfbbn_1_27/a_2136_47# 0 0.133f
C17505 sky130_fd_sc_hd__dfbbn_1_27/a_791_47# 0 0.0125f
C17506 sky130_fd_sc_hd__dfbbn_1_27/a_381_47# 0 0.0218f
C17507 sky130_fd_sc_hd__dfbbn_1_27/a_1256_413# 0 0.12f
C17508 sky130_fd_sc_hd__dfbbn_1_27/a_1415_315# 0 0.394f
C17509 sky130_fd_sc_hd__dfbbn_1_27/a_941_21# 0 0.245f
C17510 sky130_fd_sc_hd__dfbbn_1_27/a_473_413# 0 0.119f
C17511 sky130_fd_sc_hd__dfbbn_1_27/a_647_21# 0 0.24f
C17512 sky130_fd_sc_hd__dfbbn_1_27/a_193_47# 0 0.27f
C17513 sky130_fd_sc_hd__dfbbn_1_27/a_27_47# 0 0.492f
C17514 sky130_fd_sc_hd__dfbbn_1_49/Q_N 0 0.0135f
C17515 sky130_fd_sc_hd__dfbbn_1_49/a_1555_47# 0 0.00871f
C17516 sky130_fd_sc_hd__dfbbn_1_49/a_2136_47# 0 0.133f
C17517 sky130_fd_sc_hd__dfbbn_1_49/a_791_47# 0 0.0125f
C17518 sky130_fd_sc_hd__dfbbn_1_49/a_381_47# 0 0.0218f
C17519 sky130_fd_sc_hd__dfbbn_1_49/a_1256_413# 0 0.12f
C17520 sky130_fd_sc_hd__dfbbn_1_49/a_1415_315# 0 0.394f
C17521 sky130_fd_sc_hd__dfbbn_1_49/a_941_21# 0 0.245f
C17522 sky130_fd_sc_hd__dfbbn_1_49/a_473_413# 0 0.119f
C17523 sky130_fd_sc_hd__dfbbn_1_49/a_647_21# 0 0.24f
C17524 sky130_fd_sc_hd__dfbbn_1_49/a_193_47# 0 0.27f
C17525 sky130_fd_sc_hd__dfbbn_1_49/a_27_47# 0 0.492f
C17526 sky130_fd_sc_hd__dfbbn_1_38/Q_N 0 0.0135f
C17527 sky130_fd_sc_hd__dfbbn_1_38/a_1555_47# 0 0.00871f
C17528 sky130_fd_sc_hd__dfbbn_1_38/a_2136_47# 0 0.133f
C17529 sky130_fd_sc_hd__dfbbn_1_38/a_791_47# 0 0.0125f
C17530 sky130_fd_sc_hd__dfbbn_1_38/a_381_47# 0 0.0218f
C17531 sky130_fd_sc_hd__dfbbn_1_38/a_1256_413# 0 0.12f
C17532 sky130_fd_sc_hd__dfbbn_1_38/a_1415_315# 0 0.394f
C17533 sky130_fd_sc_hd__dfbbn_1_38/a_941_21# 0 0.245f
C17534 sky130_fd_sc_hd__dfbbn_1_38/a_473_413# 0 0.119f
C17535 sky130_fd_sc_hd__dfbbn_1_38/a_647_21# 0 0.24f
C17536 sky130_fd_sc_hd__dfbbn_1_38/a_193_47# 0 0.27f
C17537 sky130_fd_sc_hd__dfbbn_1_38/a_27_47# 0 0.492f
C17538 sky130_fd_sc_hd__conb_1_36/HI 0 0.474f
C17539 sky130_fd_sc_hd__inv_1_45/Y 0 0.181f
C17540 sky130_fd_sc_hd__nand2_1_2/A 0 0.165f
C17541 sky130_fd_sc_hd__conb_1_10/LO 0 0.166f
C17542 sky130_fd_sc_hd__conb_1_21/LO 0 0.166f
C17543 sky130_fd_sc_hd__conb_1_32/LO 0 0.166f
C17544 sky130_fd_sc_hd__conb_1_43/LO 0 0.166f
C17545 RISING_COUNTER.COUNT_SUB_DFF1.Q 0 0.851f
C17546 sky130_fd_sc_hd__conb_1_19/HI 0 0.464f
C17547 sky130_fd_sc_hd__dfbbn_1_26/Q_N 0 0.0135f
C17548 sky130_fd_sc_hd__dfbbn_1_26/a_1555_47# 0 0.00871f
C17549 sky130_fd_sc_hd__dfbbn_1_26/a_2136_47# 0 0.133f
C17550 sky130_fd_sc_hd__dfbbn_1_26/a_791_47# 0 0.0125f
C17551 sky130_fd_sc_hd__dfbbn_1_26/a_381_47# 0 0.0218f
C17552 sky130_fd_sc_hd__dfbbn_1_26/a_1256_413# 0 0.12f
C17553 sky130_fd_sc_hd__dfbbn_1_26/a_1415_315# 0 0.394f
C17554 sky130_fd_sc_hd__dfbbn_1_26/a_941_21# 0 0.245f
C17555 sky130_fd_sc_hd__dfbbn_1_26/a_473_413# 0 0.119f
C17556 sky130_fd_sc_hd__dfbbn_1_26/a_647_21# 0 0.24f
C17557 sky130_fd_sc_hd__dfbbn_1_26/a_193_47# 0 0.27f
C17558 sky130_fd_sc_hd__dfbbn_1_26/a_27_47# 0 0.492f
C17559 sky130_fd_sc_hd__dfbbn_1_48/Q_N 0 0.0135f
C17560 sky130_fd_sc_hd__dfbbn_1_48/a_1555_47# 0 0.00871f
C17561 sky130_fd_sc_hd__dfbbn_1_48/a_2136_47# 0 0.133f
C17562 sky130_fd_sc_hd__dfbbn_1_48/a_791_47# 0 0.0125f
C17563 sky130_fd_sc_hd__dfbbn_1_48/a_381_47# 0 0.0218f
C17564 sky130_fd_sc_hd__dfbbn_1_48/a_1256_413# 0 0.12f
C17565 sky130_fd_sc_hd__dfbbn_1_48/a_1415_315# 0 0.394f
C17566 sky130_fd_sc_hd__dfbbn_1_48/a_941_21# 0 0.245f
C17567 sky130_fd_sc_hd__dfbbn_1_48/a_473_413# 0 0.119f
C17568 sky130_fd_sc_hd__dfbbn_1_48/a_647_21# 0 0.24f
C17569 sky130_fd_sc_hd__dfbbn_1_48/a_193_47# 0 0.27f
C17570 sky130_fd_sc_hd__dfbbn_1_48/a_27_47# 0 0.492f
C17571 sky130_fd_sc_hd__dfbbn_1_37/Q_N 0 0.0135f
C17572 sky130_fd_sc_hd__dfbbn_1_37/a_1555_47# 0 0.00871f
C17573 sky130_fd_sc_hd__dfbbn_1_37/a_2136_47# 0 0.133f
C17574 sky130_fd_sc_hd__dfbbn_1_37/a_791_47# 0 0.0125f
C17575 sky130_fd_sc_hd__dfbbn_1_37/a_381_47# 0 0.0218f
C17576 sky130_fd_sc_hd__dfbbn_1_37/a_1256_413# 0 0.12f
C17577 sky130_fd_sc_hd__dfbbn_1_37/a_1415_315# 0 0.394f
C17578 sky130_fd_sc_hd__dfbbn_1_37/a_941_21# 0 0.245f
C17579 sky130_fd_sc_hd__dfbbn_1_37/a_473_413# 0 0.119f
C17580 sky130_fd_sc_hd__dfbbn_1_37/a_647_21# 0 0.24f
C17581 sky130_fd_sc_hd__dfbbn_1_37/a_193_47# 0 0.27f
C17582 sky130_fd_sc_hd__dfbbn_1_37/a_27_47# 0 0.492f
C17583 sky130_fd_sc_hd__dfbbn_1_15/Q_N 0 0.0135f
C17584 sky130_fd_sc_hd__dfbbn_1_15/a_1555_47# 0 0.00871f
C17585 sky130_fd_sc_hd__dfbbn_1_15/a_2136_47# 0 0.133f
C17586 sky130_fd_sc_hd__dfbbn_1_15/a_791_47# 0 0.0125f
C17587 sky130_fd_sc_hd__dfbbn_1_15/a_381_47# 0 0.0218f
C17588 sky130_fd_sc_hd__dfbbn_1_15/a_1256_413# 0 0.12f
C17589 sky130_fd_sc_hd__dfbbn_1_15/a_1415_315# 0 0.394f
C17590 sky130_fd_sc_hd__dfbbn_1_15/a_941_21# 0 0.245f
C17591 sky130_fd_sc_hd__dfbbn_1_15/a_473_413# 0 0.119f
C17592 sky130_fd_sc_hd__dfbbn_1_15/a_647_21# 0 0.24f
C17593 sky130_fd_sc_hd__dfbbn_1_15/a_193_47# 0 0.27f
C17594 sky130_fd_sc_hd__dfbbn_1_15/a_27_47# 0 0.492f
C17595 FALLING_COUNTER.COUNT_SUB_DFF3.Q 0 1.88f
C17596 sky130_fd_sc_hd__conb_1_20/LO 0 0.166f
C17597 sky130_fd_sc_hd__conb_1_31/LO 0 0.166f
C17598 sky130_fd_sc_hd__conb_1_42/LO 0 0.166f
C17599 sky130_fd_sc_hd__inv_1_7/Y 0 0.314f
C17600 sky130_fd_sc_hd__conb_1_10/HI 0 0.492f
C17601 sky130_fd_sc_hd__inv_1_14/Y 0 0.206f
C17602 sky130_fd_sc_hd__dfbbn_1_14/Q_N 0 0.0135f
C17603 sky130_fd_sc_hd__dfbbn_1_14/a_1555_47# 0 0.00871f
C17604 sky130_fd_sc_hd__dfbbn_1_14/a_2136_47# 0 0.133f
C17605 sky130_fd_sc_hd__dfbbn_1_14/a_791_47# 0 0.0125f
C17606 sky130_fd_sc_hd__dfbbn_1_14/a_381_47# 0 0.0218f
C17607 sky130_fd_sc_hd__dfbbn_1_14/a_1256_413# 0 0.12f
C17608 sky130_fd_sc_hd__dfbbn_1_14/a_1415_315# 0 0.394f
C17609 sky130_fd_sc_hd__dfbbn_1_14/a_941_21# 0 0.245f
C17610 sky130_fd_sc_hd__dfbbn_1_14/a_473_413# 0 0.119f
C17611 sky130_fd_sc_hd__dfbbn_1_14/a_647_21# 0 0.24f
C17612 sky130_fd_sc_hd__dfbbn_1_14/a_193_47# 0 0.27f
C17613 sky130_fd_sc_hd__dfbbn_1_14/a_27_47# 0 0.492f
C17614 sky130_fd_sc_hd__dfbbn_1_47/Q_N 0 0.0135f
C17615 sky130_fd_sc_hd__conb_1_25/HI 0 0.425f
C17616 sky130_fd_sc_hd__dfbbn_1_47/a_1555_47# 0 0.00871f
C17617 sky130_fd_sc_hd__dfbbn_1_47/a_2136_47# 0 0.133f
C17618 sky130_fd_sc_hd__dfbbn_1_47/a_791_47# 0 0.0125f
C17619 sky130_fd_sc_hd__dfbbn_1_47/a_381_47# 0 0.0218f
C17620 sky130_fd_sc_hd__dfbbn_1_47/a_1256_413# 0 0.12f
C17621 sky130_fd_sc_hd__dfbbn_1_47/a_1415_315# 0 0.394f
C17622 sky130_fd_sc_hd__dfbbn_1_47/a_941_21# 0 0.245f
C17623 sky130_fd_sc_hd__dfbbn_1_47/a_473_413# 0 0.119f
C17624 sky130_fd_sc_hd__dfbbn_1_47/a_647_21# 0 0.24f
C17625 sky130_fd_sc_hd__dfbbn_1_47/a_193_47# 0 0.27f
C17626 sky130_fd_sc_hd__dfbbn_1_47/a_27_47# 0 0.492f
C17627 sky130_fd_sc_hd__dfbbn_1_25/Q_N 0 0.0135f
C17628 sky130_fd_sc_hd__dfbbn_1_25/a_1555_47# 0 0.00871f
C17629 sky130_fd_sc_hd__dfbbn_1_25/a_2136_47# 0 0.133f
C17630 sky130_fd_sc_hd__dfbbn_1_25/a_791_47# 0 0.0125f
C17631 sky130_fd_sc_hd__dfbbn_1_25/a_381_47# 0 0.0218f
C17632 sky130_fd_sc_hd__dfbbn_1_25/a_1256_413# 0 0.12f
C17633 sky130_fd_sc_hd__dfbbn_1_25/a_1415_315# 0 0.394f
C17634 sky130_fd_sc_hd__dfbbn_1_25/a_941_21# 0 0.245f
C17635 sky130_fd_sc_hd__dfbbn_1_25/a_473_413# 0 0.119f
C17636 sky130_fd_sc_hd__dfbbn_1_25/a_647_21# 0 0.24f
C17637 sky130_fd_sc_hd__dfbbn_1_25/a_193_47# 0 0.27f
C17638 sky130_fd_sc_hd__dfbbn_1_25/a_27_47# 0 0.492f
C17639 sky130_fd_sc_hd__dfbbn_1_36/Q_N 0 0.0135f
C17640 sky130_fd_sc_hd__dfbbn_1_36/a_1555_47# 0 0.00871f
C17641 sky130_fd_sc_hd__dfbbn_1_36/a_2136_47# 0 0.133f
C17642 sky130_fd_sc_hd__dfbbn_1_36/a_791_47# 0 0.0125f
C17643 sky130_fd_sc_hd__dfbbn_1_36/a_381_47# 0 0.0218f
C17644 sky130_fd_sc_hd__dfbbn_1_36/a_1256_413# 0 0.12f
C17645 sky130_fd_sc_hd__dfbbn_1_36/a_1415_315# 0 0.394f
C17646 sky130_fd_sc_hd__dfbbn_1_36/a_941_21# 0 0.245f
C17647 sky130_fd_sc_hd__dfbbn_1_36/a_473_413# 0 0.119f
C17648 sky130_fd_sc_hd__dfbbn_1_36/a_647_21# 0 0.24f
C17649 sky130_fd_sc_hd__dfbbn_1_36/a_193_47# 0 0.27f
C17650 sky130_fd_sc_hd__dfbbn_1_36/a_27_47# 0 0.492f
C17651 sky130_fd_sc_hd__conb_1_30/LO 0 0.166f
C17652 sky130_fd_sc_hd__conb_1_41/LO 0 0.166f
C17653 sky130_fd_sc_hd__dfbbn_1_13/Q_N 0 0.0135f
C17654 sky130_fd_sc_hd__dfbbn_1_13/a_1555_47# 0 0.00871f
C17655 sky130_fd_sc_hd__dfbbn_1_13/a_2136_47# 0 0.133f
C17656 sky130_fd_sc_hd__dfbbn_1_13/a_791_47# 0 0.0125f
C17657 sky130_fd_sc_hd__dfbbn_1_13/a_381_47# 0 0.0218f
C17658 sky130_fd_sc_hd__dfbbn_1_13/a_1256_413# 0 0.12f
C17659 sky130_fd_sc_hd__dfbbn_1_13/a_1415_315# 0 0.394f
C17660 sky130_fd_sc_hd__dfbbn_1_13/a_941_21# 0 0.245f
C17661 sky130_fd_sc_hd__dfbbn_1_13/a_473_413# 0 0.119f
C17662 sky130_fd_sc_hd__dfbbn_1_13/a_647_21# 0 0.24f
C17663 sky130_fd_sc_hd__dfbbn_1_13/a_193_47# 0 0.27f
C17664 sky130_fd_sc_hd__dfbbn_1_13/a_27_47# 0 0.492f
C17665 sky130_fd_sc_hd__dfbbn_1_24/Q_N 0 0.0135f
C17666 sky130_fd_sc_hd__dfbbn_1_24/a_1555_47# 0 0.00871f
C17667 sky130_fd_sc_hd__dfbbn_1_24/a_2136_47# 0 0.133f
C17668 sky130_fd_sc_hd__dfbbn_1_24/a_791_47# 0 0.0125f
C17669 sky130_fd_sc_hd__dfbbn_1_24/a_381_47# 0 0.0218f
C17670 sky130_fd_sc_hd__dfbbn_1_24/a_1256_413# 0 0.12f
C17671 sky130_fd_sc_hd__dfbbn_1_24/a_1415_315# 0 0.394f
C17672 sky130_fd_sc_hd__dfbbn_1_24/a_941_21# 0 0.245f
C17673 sky130_fd_sc_hd__dfbbn_1_24/a_473_413# 0 0.119f
C17674 sky130_fd_sc_hd__dfbbn_1_24/a_647_21# 0 0.24f
C17675 sky130_fd_sc_hd__dfbbn_1_24/a_193_47# 0 0.27f
C17676 sky130_fd_sc_hd__dfbbn_1_24/a_27_47# 0 0.492f
C17677 sky130_fd_sc_hd__dfbbn_1_35/Q_N 0 0.0135f
C17678 sky130_fd_sc_hd__dfbbn_1_35/a_1555_47# 0 0.00871f
C17679 sky130_fd_sc_hd__dfbbn_1_35/a_2136_47# 0 0.133f
C17680 sky130_fd_sc_hd__dfbbn_1_35/a_791_47# 0 0.0125f
C17681 sky130_fd_sc_hd__dfbbn_1_35/a_381_47# 0 0.0218f
C17682 sky130_fd_sc_hd__dfbbn_1_35/a_1256_413# 0 0.12f
C17683 sky130_fd_sc_hd__dfbbn_1_35/a_1415_315# 0 0.394f
C17684 sky130_fd_sc_hd__dfbbn_1_35/a_941_21# 0 0.245f
C17685 sky130_fd_sc_hd__dfbbn_1_35/a_473_413# 0 0.119f
C17686 sky130_fd_sc_hd__dfbbn_1_35/a_647_21# 0 0.24f
C17687 sky130_fd_sc_hd__dfbbn_1_35/a_193_47# 0 0.27f
C17688 sky130_fd_sc_hd__dfbbn_1_35/a_27_47# 0 0.492f
C17689 sky130_fd_sc_hd__dfbbn_1_46/Q_N 0 0.0135f
C17690 sky130_fd_sc_hd__dfbbn_1_46/a_1555_47# 0 0.00871f
C17691 sky130_fd_sc_hd__dfbbn_1_46/a_2136_47# 0 0.133f
C17692 sky130_fd_sc_hd__dfbbn_1_46/a_791_47# 0 0.0125f
C17693 sky130_fd_sc_hd__dfbbn_1_46/a_381_47# 0 0.0218f
C17694 sky130_fd_sc_hd__dfbbn_1_46/a_1256_413# 0 0.12f
C17695 sky130_fd_sc_hd__dfbbn_1_46/a_1415_315# 0 0.394f
C17696 sky130_fd_sc_hd__dfbbn_1_46/a_941_21# 0 0.245f
C17697 sky130_fd_sc_hd__dfbbn_1_46/a_473_413# 0 0.119f
C17698 sky130_fd_sc_hd__dfbbn_1_46/a_647_21# 0 0.24f
C17699 sky130_fd_sc_hd__dfbbn_1_46/a_193_47# 0 0.27f
C17700 sky130_fd_sc_hd__dfbbn_1_46/a_27_47# 0 0.492f
C17701 sky130_fd_sc_hd__conb_1_20/HI 0 0.514f
C17702 sky130_fd_sc_hd__conb_1_51/LO 0 0.166f
C17703 sky130_fd_sc_hd__inv_1_94/Y 0 0.779f
C17704 sky130_fd_sc_hd__conb_1_40/LO 0 0.166f
C17705 sky130_fd_sc_hd__dfbbn_1_12/Q_N 0 0.0135f
C17706 sky130_fd_sc_hd__dfbbn_1_12/a_1555_47# 0 0.00871f
C17707 sky130_fd_sc_hd__dfbbn_1_12/a_2136_47# 0 0.133f
C17708 sky130_fd_sc_hd__dfbbn_1_12/a_791_47# 0 0.0125f
C17709 sky130_fd_sc_hd__dfbbn_1_12/a_381_47# 0 0.0218f
C17710 sky130_fd_sc_hd__dfbbn_1_12/a_1256_413# 0 0.12f
C17711 sky130_fd_sc_hd__dfbbn_1_12/a_1415_315# 0 0.394f
C17712 sky130_fd_sc_hd__dfbbn_1_12/a_941_21# 0 0.245f
C17713 sky130_fd_sc_hd__dfbbn_1_12/a_473_413# 0 0.119f
C17714 sky130_fd_sc_hd__dfbbn_1_12/a_647_21# 0 0.24f
C17715 sky130_fd_sc_hd__dfbbn_1_12/a_193_47# 0 0.27f
C17716 sky130_fd_sc_hd__dfbbn_1_12/a_27_47# 0 0.492f
C17717 sky130_fd_sc_hd__dfbbn_1_23/Q_N 0 0.0135f
C17718 sky130_fd_sc_hd__dfbbn_1_23/a_1555_47# 0 0.00871f
C17719 sky130_fd_sc_hd__dfbbn_1_23/a_2136_47# 0 0.133f
C17720 sky130_fd_sc_hd__dfbbn_1_23/a_791_47# 0 0.0125f
C17721 sky130_fd_sc_hd__dfbbn_1_23/a_381_47# 0 0.0218f
C17722 sky130_fd_sc_hd__dfbbn_1_23/a_1256_413# 0 0.12f
C17723 sky130_fd_sc_hd__dfbbn_1_23/a_1415_315# 0 0.394f
C17724 sky130_fd_sc_hd__dfbbn_1_23/a_941_21# 0 0.245f
C17725 sky130_fd_sc_hd__dfbbn_1_23/a_473_413# 0 0.119f
C17726 sky130_fd_sc_hd__dfbbn_1_23/a_647_21# 0 0.24f
C17727 sky130_fd_sc_hd__dfbbn_1_23/a_193_47# 0 0.27f
C17728 sky130_fd_sc_hd__dfbbn_1_23/a_27_47# 0 0.492f
C17729 sky130_fd_sc_hd__dfbbn_1_45/Q_N 0 0.0135f
C17730 sky130_fd_sc_hd__conb_1_48/HI 0 0.434f
C17731 sky130_fd_sc_hd__dfbbn_1_45/a_1555_47# 0 0.00871f
C17732 sky130_fd_sc_hd__dfbbn_1_45/a_2136_47# 0 0.133f
C17733 sky130_fd_sc_hd__dfbbn_1_45/a_791_47# 0 0.0125f
C17734 sky130_fd_sc_hd__dfbbn_1_45/a_381_47# 0 0.0218f
C17735 sky130_fd_sc_hd__dfbbn_1_45/a_1256_413# 0 0.12f
C17736 sky130_fd_sc_hd__dfbbn_1_45/a_1415_315# 0 0.394f
C17737 sky130_fd_sc_hd__dfbbn_1_45/a_941_21# 0 0.245f
C17738 sky130_fd_sc_hd__dfbbn_1_45/a_473_413# 0 0.119f
C17739 sky130_fd_sc_hd__dfbbn_1_45/a_647_21# 0 0.24f
C17740 sky130_fd_sc_hd__dfbbn_1_45/a_193_47# 0 0.27f
C17741 sky130_fd_sc_hd__dfbbn_1_45/a_27_47# 0 0.492f
C17742 sky130_fd_sc_hd__dfbbn_1_34/Q_N 0 0.0135f
C17743 sky130_fd_sc_hd__dfbbn_1_34/a_1555_47# 0 0.00871f
C17744 sky130_fd_sc_hd__dfbbn_1_34/a_2136_47# 0 0.133f
C17745 sky130_fd_sc_hd__dfbbn_1_34/a_791_47# 0 0.0125f
C17746 sky130_fd_sc_hd__dfbbn_1_34/a_381_47# 0 0.0218f
C17747 sky130_fd_sc_hd__dfbbn_1_34/a_1256_413# 0 0.12f
C17748 sky130_fd_sc_hd__dfbbn_1_34/a_1415_315# 0 0.394f
C17749 sky130_fd_sc_hd__dfbbn_1_34/a_941_21# 0 0.245f
C17750 sky130_fd_sc_hd__dfbbn_1_34/a_473_413# 0 0.119f
C17751 sky130_fd_sc_hd__dfbbn_1_34/a_647_21# 0 0.24f
C17752 sky130_fd_sc_hd__dfbbn_1_34/a_193_47# 0 0.27f
C17753 sky130_fd_sc_hd__dfbbn_1_34/a_27_47# 0 0.492f
C17754 sky130_fd_sc_hd__conb_1_50/LO 0 0.166f
C17755 sky130_fd_sc_hd__inv_1_96/A 0 0.436f
C17756 sky130_fd_sc_hd__dfbbn_1_44/Q_N 0 0.0135f
C17757 sky130_fd_sc_hd__dfbbn_1_44/a_1555_47# 0 0.00871f
C17758 sky130_fd_sc_hd__dfbbn_1_44/a_2136_47# 0 0.133f
C17759 sky130_fd_sc_hd__dfbbn_1_44/a_791_47# 0 0.0125f
C17760 sky130_fd_sc_hd__dfbbn_1_44/a_381_47# 0 0.0218f
C17761 sky130_fd_sc_hd__dfbbn_1_44/a_1256_413# 0 0.12f
C17762 sky130_fd_sc_hd__dfbbn_1_44/a_1415_315# 0 0.394f
C17763 sky130_fd_sc_hd__dfbbn_1_44/a_941_21# 0 0.245f
C17764 sky130_fd_sc_hd__dfbbn_1_44/a_473_413# 0 0.119f
C17765 sky130_fd_sc_hd__dfbbn_1_44/a_647_21# 0 0.24f
C17766 sky130_fd_sc_hd__dfbbn_1_44/a_193_47# 0 0.27f
C17767 sky130_fd_sc_hd__dfbbn_1_44/a_27_47# 0 0.492f
C17768 sky130_fd_sc_hd__dfbbn_1_11/Q_N 0 0.0135f
C17769 sky130_fd_sc_hd__dfbbn_1_11/a_1555_47# 0 0.00871f
C17770 sky130_fd_sc_hd__dfbbn_1_11/a_2136_47# 0 0.133f
C17771 sky130_fd_sc_hd__dfbbn_1_11/a_791_47# 0 0.0125f
C17772 sky130_fd_sc_hd__dfbbn_1_11/a_381_47# 0 0.0218f
C17773 sky130_fd_sc_hd__dfbbn_1_11/a_1256_413# 0 0.12f
C17774 sky130_fd_sc_hd__dfbbn_1_11/a_1415_315# 0 0.394f
C17775 sky130_fd_sc_hd__dfbbn_1_11/a_941_21# 0 0.245f
C17776 sky130_fd_sc_hd__dfbbn_1_11/a_473_413# 0 0.119f
C17777 sky130_fd_sc_hd__dfbbn_1_11/a_647_21# 0 0.24f
C17778 sky130_fd_sc_hd__dfbbn_1_11/a_193_47# 0 0.27f
C17779 sky130_fd_sc_hd__dfbbn_1_11/a_27_47# 0 0.492f
C17780 sky130_fd_sc_hd__dfbbn_1_22/Q_N 0 0.0135f
C17781 sky130_fd_sc_hd__dfbbn_1_22/a_1555_47# 0 0.00871f
C17782 sky130_fd_sc_hd__dfbbn_1_22/a_2136_47# 0 0.133f
C17783 sky130_fd_sc_hd__dfbbn_1_22/a_791_47# 0 0.0125f
C17784 sky130_fd_sc_hd__dfbbn_1_22/a_381_47# 0 0.0218f
C17785 sky130_fd_sc_hd__dfbbn_1_22/a_1256_413# 0 0.12f
C17786 sky130_fd_sc_hd__dfbbn_1_22/a_1415_315# 0 0.394f
C17787 sky130_fd_sc_hd__dfbbn_1_22/a_941_21# 0 0.245f
C17788 sky130_fd_sc_hd__dfbbn_1_22/a_473_413# 0 0.119f
C17789 sky130_fd_sc_hd__dfbbn_1_22/a_647_21# 0 0.24f
C17790 sky130_fd_sc_hd__dfbbn_1_22/a_193_47# 0 0.27f
C17791 sky130_fd_sc_hd__dfbbn_1_22/a_27_47# 0 0.492f
C17792 sky130_fd_sc_hd__dfbbn_1_33/Q_N 0 0.0135f
C17793 sky130_fd_sc_hd__dfbbn_1_33/a_1555_47# 0 0.00871f
C17794 sky130_fd_sc_hd__dfbbn_1_33/a_2136_47# 0 0.133f
C17795 sky130_fd_sc_hd__dfbbn_1_33/a_791_47# 0 0.0125f
C17796 sky130_fd_sc_hd__dfbbn_1_33/a_381_47# 0 0.0218f
C17797 sky130_fd_sc_hd__dfbbn_1_33/a_1256_413# 0 0.12f
C17798 sky130_fd_sc_hd__dfbbn_1_33/a_1415_315# 0 0.394f
C17799 sky130_fd_sc_hd__dfbbn_1_33/a_941_21# 0 0.245f
C17800 sky130_fd_sc_hd__dfbbn_1_33/a_473_413# 0 0.119f
C17801 sky130_fd_sc_hd__dfbbn_1_33/a_647_21# 0 0.24f
C17802 sky130_fd_sc_hd__dfbbn_1_33/a_193_47# 0 0.27f
C17803 sky130_fd_sc_hd__dfbbn_1_33/a_27_47# 0 0.492f
C17804 FALLING_COUNTER.COUNT_SUB_DFF6.Q 0 1.87f
C17805 sky130_fd_sc_hd__inv_1_110/Y 0 0.264f
C17806 sky130_fd_sc_hd__dfbbn_1_10/Q_N 0 0.0135f
C17807 sky130_fd_sc_hd__dfbbn_1_10/a_1555_47# 0 0.00871f
C17808 sky130_fd_sc_hd__dfbbn_1_10/a_2136_47# 0 0.133f
C17809 sky130_fd_sc_hd__dfbbn_1_10/a_791_47# 0 0.0125f
C17810 sky130_fd_sc_hd__dfbbn_1_10/a_381_47# 0 0.0218f
C17811 sky130_fd_sc_hd__dfbbn_1_10/a_1256_413# 0 0.12f
C17812 sky130_fd_sc_hd__dfbbn_1_10/a_1415_315# 0 0.394f
C17813 sky130_fd_sc_hd__dfbbn_1_10/a_941_21# 0 0.245f
C17814 sky130_fd_sc_hd__dfbbn_1_10/a_473_413# 0 0.119f
C17815 sky130_fd_sc_hd__dfbbn_1_10/a_647_21# 0 0.24f
C17816 sky130_fd_sc_hd__dfbbn_1_10/a_193_47# 0 0.27f
C17817 sky130_fd_sc_hd__dfbbn_1_10/a_27_47# 0 0.492f
C17818 sky130_fd_sc_hd__dfbbn_1_21/Q_N 0 0.0135f
C17819 sky130_fd_sc_hd__dfbbn_1_21/a_1555_47# 0 0.00871f
C17820 sky130_fd_sc_hd__dfbbn_1_21/a_2136_47# 0 0.133f
C17821 sky130_fd_sc_hd__dfbbn_1_21/a_791_47# 0 0.0125f
C17822 sky130_fd_sc_hd__dfbbn_1_21/a_381_47# 0 0.0218f
C17823 sky130_fd_sc_hd__dfbbn_1_21/a_1256_413# 0 0.12f
C17824 sky130_fd_sc_hd__dfbbn_1_21/a_1415_315# 0 0.394f
C17825 sky130_fd_sc_hd__dfbbn_1_21/a_941_21# 0 0.245f
C17826 sky130_fd_sc_hd__dfbbn_1_21/a_473_413# 0 0.119f
C17827 sky130_fd_sc_hd__dfbbn_1_21/a_647_21# 0 0.24f
C17828 sky130_fd_sc_hd__dfbbn_1_21/a_193_47# 0 0.27f
C17829 sky130_fd_sc_hd__dfbbn_1_21/a_27_47# 0 0.492f
C17830 sky130_fd_sc_hd__dfbbn_1_43/Q_N 0 0.0135f
C17831 sky130_fd_sc_hd__dfbbn_1_43/a_1555_47# 0 0.00871f
C17832 sky130_fd_sc_hd__dfbbn_1_43/a_2136_47# 0 0.133f
C17833 sky130_fd_sc_hd__dfbbn_1_43/a_791_47# 0 0.0125f
C17834 sky130_fd_sc_hd__dfbbn_1_43/a_381_47# 0 0.0218f
C17835 sky130_fd_sc_hd__dfbbn_1_43/a_1256_413# 0 0.12f
C17836 sky130_fd_sc_hd__dfbbn_1_43/a_1415_315# 0 0.394f
C17837 sky130_fd_sc_hd__dfbbn_1_43/a_941_21# 0 0.245f
C17838 sky130_fd_sc_hd__dfbbn_1_43/a_473_413# 0 0.119f
C17839 sky130_fd_sc_hd__dfbbn_1_43/a_647_21# 0 0.24f
C17840 sky130_fd_sc_hd__dfbbn_1_43/a_193_47# 0 0.27f
C17841 sky130_fd_sc_hd__dfbbn_1_43/a_27_47# 0 0.492f
C17842 sky130_fd_sc_hd__dfbbn_1_32/Q_N 0 0.0135f
C17843 sky130_fd_sc_hd__dfbbn_1_32/a_1555_47# 0 0.00871f
C17844 sky130_fd_sc_hd__dfbbn_1_32/a_2136_47# 0 0.133f
C17845 sky130_fd_sc_hd__dfbbn_1_32/a_791_47# 0 0.0125f
C17846 sky130_fd_sc_hd__dfbbn_1_32/a_381_47# 0 0.0218f
C17847 sky130_fd_sc_hd__dfbbn_1_32/a_1256_413# 0 0.12f
C17848 sky130_fd_sc_hd__dfbbn_1_32/a_1415_315# 0 0.394f
C17849 sky130_fd_sc_hd__dfbbn_1_32/a_941_21# 0 0.245f
C17850 sky130_fd_sc_hd__dfbbn_1_32/a_473_413# 0 0.119f
C17851 sky130_fd_sc_hd__dfbbn_1_32/a_647_21# 0 0.24f
C17852 sky130_fd_sc_hd__dfbbn_1_32/a_193_47# 0 0.27f
C17853 sky130_fd_sc_hd__dfbbn_1_32/a_27_47# 0 0.492f
C17854 FALLING_COUNTER.COUNT_SUB_DFF4.Q 0 1.6f
C17855 sky130_fd_sc_hd__inv_1_104/Y 0 0.174f
C17856 sky130_fd_sc_hd__inv_1_17/Y 0 0.194f
C17857 sky130_fd_sc_hd__inv_1_46/A 0 0.258f
C17858 sky130_fd_sc_hd__inv_1_96/Y 0 0.681f
C17859 sky130_fd_sc_hd__inv_1_64/Y 0 0.13f
C17860 sky130_fd_sc_hd__conb_1_1/HI 0 0.474f
C17861 sky130_fd_sc_hd__dfbbn_1_20/Q_N 0 0.0135f
C17862 sky130_fd_sc_hd__dfbbn_1_20/a_1555_47# 0 0.00871f
C17863 sky130_fd_sc_hd__dfbbn_1_20/a_2136_47# 0 0.133f
C17864 sky130_fd_sc_hd__dfbbn_1_20/a_791_47# 0 0.0125f
C17865 sky130_fd_sc_hd__dfbbn_1_20/a_381_47# 0 0.0218f
C17866 sky130_fd_sc_hd__dfbbn_1_20/a_1256_413# 0 0.12f
C17867 sky130_fd_sc_hd__dfbbn_1_20/a_1415_315# 0 0.394f
C17868 sky130_fd_sc_hd__dfbbn_1_20/a_941_21# 0 0.245f
C17869 sky130_fd_sc_hd__dfbbn_1_20/a_473_413# 0 0.119f
C17870 sky130_fd_sc_hd__dfbbn_1_20/a_647_21# 0 0.24f
C17871 sky130_fd_sc_hd__dfbbn_1_20/a_193_47# 0 0.27f
C17872 sky130_fd_sc_hd__dfbbn_1_20/a_27_47# 0 0.492f
C17873 sky130_fd_sc_hd__dfbbn_1_42/Q_N 0 0.0135f
C17874 sky130_fd_sc_hd__dfbbn_1_42/a_1555_47# 0 0.00871f
C17875 sky130_fd_sc_hd__dfbbn_1_42/a_2136_47# 0 0.133f
C17876 sky130_fd_sc_hd__dfbbn_1_42/a_791_47# 0 0.0125f
C17877 sky130_fd_sc_hd__dfbbn_1_42/a_381_47# 0 0.0218f
C17878 sky130_fd_sc_hd__dfbbn_1_42/a_1256_413# 0 0.12f
C17879 sky130_fd_sc_hd__dfbbn_1_42/a_1415_315# 0 0.394f
C17880 sky130_fd_sc_hd__dfbbn_1_42/a_941_21# 0 0.245f
C17881 sky130_fd_sc_hd__dfbbn_1_42/a_473_413# 0 0.119f
C17882 sky130_fd_sc_hd__dfbbn_1_42/a_647_21# 0 0.24f
C17883 sky130_fd_sc_hd__dfbbn_1_42/a_193_47# 0 0.27f
C17884 sky130_fd_sc_hd__dfbbn_1_42/a_27_47# 0 0.492f
C17885 sky130_fd_sc_hd__dfbbn_1_31/Q_N 0 0.0135f
C17886 sky130_fd_sc_hd__dfbbn_1_31/a_1555_47# 0 0.00871f
C17887 sky130_fd_sc_hd__dfbbn_1_31/a_2136_47# 0 0.133f
C17888 sky130_fd_sc_hd__dfbbn_1_31/a_791_47# 0 0.0125f
C17889 sky130_fd_sc_hd__dfbbn_1_31/a_381_47# 0 0.0218f
C17890 sky130_fd_sc_hd__dfbbn_1_31/a_1256_413# 0 0.12f
C17891 sky130_fd_sc_hd__dfbbn_1_31/a_1415_315# 0 0.394f
C17892 sky130_fd_sc_hd__dfbbn_1_31/a_941_21# 0 0.245f
C17893 sky130_fd_sc_hd__dfbbn_1_31/a_473_413# 0 0.119f
C17894 sky130_fd_sc_hd__dfbbn_1_31/a_647_21# 0 0.24f
C17895 sky130_fd_sc_hd__dfbbn_1_31/a_193_47# 0 0.27f
C17896 sky130_fd_sc_hd__dfbbn_1_31/a_27_47# 0 0.492f
C17897 sky130_fd_sc_hd__fill_4_75/VPB 0 4.66f
C17898 sky130_fd_sc_hd__dfbbn_1_41/Q_N 0 0.0135f
C17899 sky130_fd_sc_hd__dfbbn_1_41/a_1555_47# 0 0.00871f
C17900 sky130_fd_sc_hd__dfbbn_1_41/a_2136_47# 0 0.133f
C17901 sky130_fd_sc_hd__dfbbn_1_41/a_791_47# 0 0.0125f
C17902 sky130_fd_sc_hd__dfbbn_1_41/a_381_47# 0 0.0218f
C17903 sky130_fd_sc_hd__dfbbn_1_41/a_1256_413# 0 0.12f
C17904 sky130_fd_sc_hd__dfbbn_1_41/a_1415_315# 0 0.394f
C17905 sky130_fd_sc_hd__dfbbn_1_41/a_941_21# 0 0.245f
C17906 sky130_fd_sc_hd__dfbbn_1_41/a_473_413# 0 0.119f
C17907 sky130_fd_sc_hd__dfbbn_1_41/a_647_21# 0 0.24f
C17908 sky130_fd_sc_hd__dfbbn_1_41/a_193_47# 0 0.27f
C17909 sky130_fd_sc_hd__dfbbn_1_41/a_27_47# 0 0.492f
C17910 sky130_fd_sc_hd__dfbbn_1_30/Q_N 0 0.0135f
C17911 sky130_fd_sc_hd__dfbbn_1_30/a_1555_47# 0 0.00871f
C17912 sky130_fd_sc_hd__dfbbn_1_30/a_2136_47# 0 0.133f
C17913 sky130_fd_sc_hd__dfbbn_1_30/a_791_47# 0 0.0125f
C17914 sky130_fd_sc_hd__dfbbn_1_30/a_381_47# 0 0.0218f
C17915 sky130_fd_sc_hd__dfbbn_1_30/a_1256_413# 0 0.12f
C17916 sky130_fd_sc_hd__dfbbn_1_30/a_1415_315# 0 0.394f
C17917 sky130_fd_sc_hd__dfbbn_1_30/a_941_21# 0 0.245f
C17918 sky130_fd_sc_hd__dfbbn_1_30/a_473_413# 0 0.119f
C17919 sky130_fd_sc_hd__dfbbn_1_30/a_647_21# 0 0.24f
C17920 sky130_fd_sc_hd__dfbbn_1_30/a_193_47# 0 0.27f
C17921 sky130_fd_sc_hd__dfbbn_1_30/a_27_47# 0 0.492f
C17922 sky130_fd_sc_hd__conb_1_43/HI 0 0.454f
C17923 sky130_fd_sc_hd__fill_4_74/VPB 0 4.66f
C17924 sky130_fd_sc_hd__dfbbn_1_51/Q_N 0 0.0135f
C17925 sky130_fd_sc_hd__dfbbn_1_51/a_1555_47# 0 0.00871f
C17926 sky130_fd_sc_hd__dfbbn_1_51/a_2136_47# 0 0.133f
C17927 sky130_fd_sc_hd__dfbbn_1_51/a_791_47# 0 0.0125f
C17928 sky130_fd_sc_hd__dfbbn_1_51/a_381_47# 0 0.0218f
C17929 sky130_fd_sc_hd__dfbbn_1_51/a_1256_413# 0 0.12f
C17930 sky130_fd_sc_hd__dfbbn_1_51/a_1415_315# 0 0.394f
C17931 sky130_fd_sc_hd__dfbbn_1_51/a_941_21# 0 0.245f
C17932 sky130_fd_sc_hd__dfbbn_1_51/a_473_413# 0 0.119f
C17933 sky130_fd_sc_hd__dfbbn_1_51/a_647_21# 0 0.24f
C17934 sky130_fd_sc_hd__dfbbn_1_51/a_193_47# 0 0.27f
C17935 sky130_fd_sc_hd__dfbbn_1_51/a_27_47# 0 0.492f
C17936 sky130_fd_sc_hd__dfbbn_1_40/Q_N 0 0.0135f
C17937 sky130_fd_sc_hd__dfbbn_1_40/a_1555_47# 0 0.00871f
C17938 sky130_fd_sc_hd__dfbbn_1_40/a_2136_47# 0 0.133f
C17939 sky130_fd_sc_hd__dfbbn_1_40/a_791_47# 0 0.0125f
C17940 sky130_fd_sc_hd__dfbbn_1_40/a_381_47# 0 0.0218f
C17941 sky130_fd_sc_hd__dfbbn_1_40/a_1256_413# 0 0.12f
C17942 sky130_fd_sc_hd__dfbbn_1_40/a_1415_315# 0 0.394f
C17943 sky130_fd_sc_hd__dfbbn_1_40/a_941_21# 0 0.245f
C17944 sky130_fd_sc_hd__dfbbn_1_40/a_473_413# 0 0.119f
C17945 sky130_fd_sc_hd__dfbbn_1_40/a_647_21# 0 0.24f
C17946 sky130_fd_sc_hd__dfbbn_1_40/a_193_47# 0 0.27f
C17947 sky130_fd_sc_hd__dfbbn_1_40/a_27_47# 0 0.492f
C17948 sky130_fd_sc_hd__inv_1_49/Y 0 0.296f
C17949 sky130_fd_sc_hd__fill_4_69/VPB 0 4.66f
C17950 sky130_fd_sc_hd__dfbbn_1_50/Q_N 0 0.0135f
C17951 sky130_fd_sc_hd__dfbbn_1_50/a_1555_47# 0 0.00871f
C17952 sky130_fd_sc_hd__dfbbn_1_50/a_2136_47# 0 0.133f
C17953 sky130_fd_sc_hd__dfbbn_1_50/a_791_47# 0 0.0125f
C17954 sky130_fd_sc_hd__dfbbn_1_50/a_381_47# 0 0.0218f
C17955 sky130_fd_sc_hd__dfbbn_1_50/a_1256_413# 0 0.12f
C17956 sky130_fd_sc_hd__dfbbn_1_50/a_1415_315# 0 0.394f
C17957 sky130_fd_sc_hd__dfbbn_1_50/a_941_21# 0 0.245f
C17958 sky130_fd_sc_hd__dfbbn_1_50/a_473_413# 0 0.119f
C17959 sky130_fd_sc_hd__dfbbn_1_50/a_647_21# 0 0.24f
C17960 sky130_fd_sc_hd__dfbbn_1_50/a_193_47# 0 0.27f
C17961 sky130_fd_sc_hd__dfbbn_1_50/a_27_47# 0 0.492f
C17962 sky130_fd_sc_hd__conb_1_7/HI 0 0.503f
C17963 sky130_fd_sc_hd__fill_4_56/VPB 0 4.66f
C17964 FALLING_COUNTER.COUNT_SUB_DFF14.Q 0 0.938f
C17965 sky130_fd_sc_hd__inv_1_89/Y 0 0.176f
C17966 sky130_fd_sc_hd__conb_1_15/HI 0 0.492f
C17967 RISING_COUNTER.COUNT_SUB_DFF14.Q 0 0.78f
C17968 sky130_fd_sc_hd__inv_1_52/Y 0 0.234f
C17969 sky130_fd_sc_hd__nand2_8_3/A 0 0.668f
C17970 sky130_fd_sc_hd__inv_1_89/A 0 0.164f
C17971 sky130_fd_sc_hd__conb_1_50/HI 0 0.468f
C17972 sky130_fd_sc_hd__nand2_8_9/a_27_47# 0 0.083f
C17973 sky130_fd_sc_hd__fill_4_58/VPB 0 4.66f
C17974 sky130_fd_sc_hd__nand2_1_5/Y 0 0.188f
C17975 sky130_fd_sc_hd__fill_4_85/VPB 0 4.66f
C17976 sky130_fd_sc_hd__nand2_8_8/a_27_47# 0 0.083f
C17977 FULL_COUNTER.COUNT_SUB_DFF12.Q 0 1.04f
C17978 sky130_fd_sc_hd__inv_1_39/Y 0 0.183f
C17979 sky130_fd_sc_hd__inv_1_48/Y 0 0.16f
C17980 sky130_fd_sc_hd__fill_4_68/VPB 0 4.66f
C17981 sky130_fd_sc_hd__fill_4_87/VPB 0 4.66f
C17982 sky130_fd_sc_hd__nand2_8_7/a_27_47# 0 0.083f
C17983 FULL_COUNTER.COUNT_SUB_DFF0.Q 0 -1.59f
C17984 sky130_fd_sc_hd__nand2_8_6/a_27_47# 0 0.083f
C17985 FULL_COUNTER.COUNT_SUB_DFF17.Q 0 1.16f
C17986 sky130_fd_sc_hd__inv_1_46/Y 0 0.212f
C17987 sky130_fd_sc_hd__inv_1_111/Y 0 0.213f
C17988 sky130_fd_sc_hd__fill_4_60/VPB 0 4.66f
C17989 sky130_fd_sc_hd__conb_1_29/HI 0 0.461f
C17990 sky130_fd_sc_hd__dfbbn_1_9/Q_N 0 0.0135f
C17991 sky130_fd_sc_hd__dfbbn_1_9/a_1555_47# 0 0.00871f
C17992 sky130_fd_sc_hd__dfbbn_1_9/a_2136_47# 0 0.133f
C17993 sky130_fd_sc_hd__dfbbn_1_9/a_791_47# 0 0.0125f
C17994 sky130_fd_sc_hd__dfbbn_1_9/a_381_47# 0 0.0218f
C17995 sky130_fd_sc_hd__dfbbn_1_9/a_1256_413# 0 0.12f
C17996 sky130_fd_sc_hd__dfbbn_1_9/a_1415_315# 0 0.394f
C17997 sky130_fd_sc_hd__dfbbn_1_9/a_941_21# 0 0.245f
C17998 sky130_fd_sc_hd__dfbbn_1_9/a_473_413# 0 0.119f
C17999 sky130_fd_sc_hd__dfbbn_1_9/a_647_21# 0 0.24f
C18000 sky130_fd_sc_hd__dfbbn_1_9/a_193_47# 0 0.27f
C18001 sky130_fd_sc_hd__dfbbn_1_9/a_27_47# 0 0.492f
C18002 sky130_fd_sc_hd__nand2_8_5/a_27_47# 0 0.083f
C18003 FULL_COUNTER.COUNT_SUB_DFF15.Q 0 1.07f
C18004 FULL_COUNTER.COUNT_SUB_DFF6.Q 0 0.993f
C18005 RISING_COUNTER.COUNT_SUB_DFF8.Q 0 0.974f
C18006 sky130_fd_sc_hd__fill_4_72/VPB 0 4.66f
C18007 sky130_fd_sc_hd__dfbbn_1_8/Q_N 0 0.0135f
C18008 sky130_fd_sc_hd__dfbbn_1_8/a_1555_47# 0 0.00871f
C18009 sky130_fd_sc_hd__dfbbn_1_8/a_2136_47# 0 0.133f
C18010 sky130_fd_sc_hd__dfbbn_1_8/a_791_47# 0 0.0125f
C18011 sky130_fd_sc_hd__dfbbn_1_8/a_381_47# 0 0.0218f
C18012 sky130_fd_sc_hd__dfbbn_1_8/a_1256_413# 0 0.12f
C18013 sky130_fd_sc_hd__dfbbn_1_8/a_1415_315# 0 0.394f
C18014 sky130_fd_sc_hd__dfbbn_1_8/a_941_21# 0 0.245f
C18015 sky130_fd_sc_hd__dfbbn_1_8/a_473_413# 0 0.119f
C18016 sky130_fd_sc_hd__dfbbn_1_8/a_647_21# 0 0.24f
C18017 sky130_fd_sc_hd__dfbbn_1_8/a_193_47# 0 0.27f
C18018 sky130_fd_sc_hd__dfbbn_1_8/a_27_47# 0 0.492f
C18019 sky130_fd_sc_hd__nand2_8_4/a_27_47# 0 0.083f
C18020 sky130_fd_sc_hd__conb_1_14/HI 0 0.509f
C18021 FALLING_COUNTER.COUNT_SUB_DFF15.Q 0 0.925f
C18022 FALLING_COUNTER.COUNT_SUB_DFF2.Q 0 1.58f
C18023 sky130_fd_sc_hd__fill_4_63/VPB 0 4.66f
C18024 sky130_fd_sc_hd__inv_1_81/Y 0 0.755f
C18025 sky130_fd_sc_hd__dfbbn_1_7/Q_N 0 0.0135f
C18026 sky130_fd_sc_hd__dfbbn_1_7/a_1555_47# 0 0.00871f
C18027 sky130_fd_sc_hd__dfbbn_1_7/a_2136_47# 0 0.133f
C18028 sky130_fd_sc_hd__dfbbn_1_7/a_791_47# 0 0.0125f
C18029 sky130_fd_sc_hd__dfbbn_1_7/a_381_47# 0 0.0218f
C18030 sky130_fd_sc_hd__dfbbn_1_7/a_1256_413# 0 0.12f
C18031 sky130_fd_sc_hd__dfbbn_1_7/a_1415_315# 0 0.394f
C18032 sky130_fd_sc_hd__dfbbn_1_7/a_941_21# 0 0.245f
C18033 sky130_fd_sc_hd__dfbbn_1_7/a_473_413# 0 0.119f
C18034 sky130_fd_sc_hd__dfbbn_1_7/a_647_21# 0 0.24f
C18035 sky130_fd_sc_hd__dfbbn_1_7/a_193_47# 0 0.27f
C18036 sky130_fd_sc_hd__dfbbn_1_7/a_27_47# 0 0.492f
C18037 sky130_fd_sc_hd__nand2_8_3/a_27_47# 0 0.083f
C18038 sky130_fd_sc_hd__fill_8_819/VPB 0 4.66f
C18039 sky130_fd_sc_hd__dfbbn_1_6/Q_N 0 0.0135f
C18040 sky130_fd_sc_hd__dfbbn_1_6/a_1555_47# 0 0.00871f
C18041 sky130_fd_sc_hd__dfbbn_1_6/a_2136_47# 0 0.133f
C18042 sky130_fd_sc_hd__dfbbn_1_6/a_791_47# 0 0.0125f
C18043 sky130_fd_sc_hd__dfbbn_1_6/a_381_47# 0 0.0218f
C18044 sky130_fd_sc_hd__dfbbn_1_6/a_1256_413# 0 0.12f
C18045 sky130_fd_sc_hd__dfbbn_1_6/a_1415_315# 0 0.394f
C18046 sky130_fd_sc_hd__dfbbn_1_6/a_941_21# 0 0.245f
C18047 sky130_fd_sc_hd__dfbbn_1_6/a_473_413# 0 0.119f
C18048 sky130_fd_sc_hd__dfbbn_1_6/a_647_21# 0 0.24f
C18049 sky130_fd_sc_hd__dfbbn_1_6/a_193_47# 0 0.27f
C18050 sky130_fd_sc_hd__dfbbn_1_6/a_27_47# 0 0.492f
C18051 sky130_fd_sc_hd__nand2_8_2/a_27_47# 0 0.083f
C18052 FULL_COUNTER.COUNT_SUB_DFF19.Q 0 1.15f
C18053 FULL_COUNTER.COUNT_SUB_DFF14.Q 0 1.41f
.ends

